------------------------------------------HEADER START"------------------------------------------
--THIS FILE WAS GENERATED USING HIGH LANGUAGE DESCRIPTION TOOL DESIGNED BY: MUHAMMAD HAMDAN
--TOOL VERSION: 0.1
--GENERATION DATE/TIME:Mon Apr 06 11:20:12 CDT 2020
------------------------------------------HEADER END"--------------------------------------------



------------------------------DESCRIPTION AND LIBRARY DECLARATION-START---------------------------
-- Engineer:       Muhammad Hamdan
-- Design Name:    HDL GENERATION - CONV LAYER 
-- Module Name:    FC - Behavioral 
-- Project Name:   CNN accelerator
-- Number of Total Operaiton: 40
-- Number of Clock Cycles: 58
-- Number of GOPS = 0.0
-------------------------------------------------Total Number of Operations for the Entire Model:10
-- Target Devices: Zynq-XC7Z020
-- Description: 
-- Dependencies: 
-- Revision:0.010 


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_arith.all;

entity FC_LAYER_8 is

GENERIC
 	( 
	constant PERCISION      : positive := 5; 	
	constant DOUT_WIDTH     : positive := 5; 	
	constant BIAS_SIZE      : positive := 5;
	constant MULT_SIZE      : positive := 10;
	constant BASE_DIN_WIDTH : positive := 75;
	constant DIN_WIDTH      : positive := 5;
	constant IMAGE_WIDTH    : positive := 1;
	constant IMAGE_SIZE     : positive := 1024;	
	constant F_SIZE         : positive := 1;
	constant PF_X2_SIZE     : positive := 25;
	constant WEIGHT_SIZE    : positive := 5;
	constant BIASES_SIZE	: positive := 2;
	constant PADDING        : positive := 1;
	constant STRIDE         : positive := 1;
	constant FEATURE_MAPS   : positive := 10;
	constant VALID_CYCLES   : positive := 25;
	constant VALID_LOCAL_PIX: positive := 5;
	constant ADD_TREE_DEPTH : positive := 1;
	constant INPUT_DEPTH    : positive := 7;
	constant INNER_PXL_SUM  : positive := 1;
	constant SUM_PEXILS     : positive := 100;
	constant MULT_SUM_D_1   : positive := 42;
	constant MULT_SUM_SIZE_1: positive := 6;
	constant MULT_SUM_D_2   : positive := 21;
	constant MULT_SUM_SIZE_2: positive := 6;
	constant MULT_SUM_D_3   : positive := 11;
	constant MULT_SUM_SIZE_3: positive := 6;
	constant MULT_SUM_D_4   : positive := 6;
	constant MULT_SUM_SIZE_4: positive := 6;
	constant MULT_SUM_D_5   : positive := 3;
	constant MULT_SUM_SIZE_5: positive := 6;
	constant MULT_SUM_D_6   : positive := 2;
	constant MULT_SUM_SIZE_6: positive := 6;
	constant MULT_SUM_D_7   : positive := 1;
	constant MULT_SUM_SIZE_7: positive := 6;
	constant LOCAL_OUTPUT   : positive := 5	
		); 

port(
	DIN_1_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_2_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_3_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_4_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_5_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_6_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_7_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_8_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_9_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_10_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_11_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_12_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_13_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_14_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_15_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_16_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_17_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_18_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_19_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_20_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_21_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_22_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_23_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_24_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_25_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_26_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_27_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_28_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_29_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_30_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_31_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_32_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_33_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_34_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_35_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_36_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_37_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_38_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_39_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_40_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_41_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_42_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_43_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_44_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_45_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_46_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_47_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_48_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_49_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_50_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_51_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_52_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_53_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_54_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_55_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_56_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_57_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_58_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_59_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_60_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_61_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_62_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_63_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_64_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_65_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_66_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_67_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_68_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_69_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_70_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_71_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_72_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_73_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_74_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_75_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_76_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_77_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_78_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_79_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_80_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_81_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_82_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_83_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_84_8         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	CLK,RST         :IN std_logic;
   	DIS_STREAM      :OUT std_logic; 				-- S_AXIS_TVALID  : Data in is valid
   	EN_STREAM       :IN std_logic; 					-- S_AXIS_TREADY  : Ready to accept data in 
	EN_STREAM_OUT_8 :OUT std_logic; 			-- M_AXIS_TREADY  : Connected slave device is ready to accept data out/ Internal Enable
	VALID_OUT_8     :OUT std_logic;                         -- M_AXIS_TVALID  : Data out is valid
	EN_LOC_STREAM_8 :IN std_logic;
	DOUT_1_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_2_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_3_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_4_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_5_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_6_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_7_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_8_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_9_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_10_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	INTERNAL_RST    :OUT std_logic
	);	

end FC_LAYER_8;

------------------------------ ARCHITECTURE DECLARATION - START---------------------------------------------

architecture Behavioral of FC_LAYER_8 is

------------------------------ INTERNAL FIXED CONSTANT & SIGNALS DECLARATION - START---------------------------------------------
type       FILTER_TYPE             is array (0 to PF_X2_SIZE-1) of signed(WEIGHT_SIZE- 1 downto 0);
signal     VALID_NXTLYR_PIX        :integer range 0 to VALID_CYCLES;
signal     PIXEL_COUNT             :integer range 0 to VALID_CYCLES;
signal     OUT_PIXEL_COUNT         :integer range 0 to VALID_CYCLES;
signal     EN_NXT_LYR_8            :std_logic;
signal     FRST_TIM_EN_8           :std_logic;
signal     Enable_MULT             :std_logic;
signal     Enable_ADDER            :std_logic;
signal     Enable_ReLU             :std_logic;
signal     Enable_BIAS             :std_logic;
signal     COUNT_PIX               :integer range 0 to PF_X2_SIZE;
signal     SIG_STRIDE              :integer range 0 to IMAGE_SIZE;
signal     PADDING_count           :integer range 0 to IMAGE_SIZE; -- TEMPORARY
signal     ROW_COUNT               :integer range 0 to IMAGE_SIZE; -- TEMPORARY


------------------------------ INTERNAL DYNAMIC SIGNALS DECLARATION ARRAY TYPE- START---------------------------------------------


type   MULT_X		is array (0 to FEATURE_MAPS-1) of signed(MULT_SIZE- 1 downto 0);
signal MULT_1:MULT_X;
signal MULT_2:MULT_X;
signal MULT_3:MULT_X;
signal MULT_4:MULT_X;
signal MULT_5:MULT_X;
signal MULT_6:MULT_X;
signal MULT_7:MULT_X;
signal MULT_8:MULT_X;
signal MULT_9:MULT_X;
signal MULT_10:MULT_X;
signal MULT_11:MULT_X;
signal MULT_12:MULT_X;
signal MULT_13:MULT_X;
signal MULT_14:MULT_X;
signal MULT_15:MULT_X;
signal MULT_16:MULT_X;
signal MULT_17:MULT_X;
signal MULT_18:MULT_X;
signal MULT_19:MULT_X;
signal MULT_20:MULT_X;
signal MULT_21:MULT_X;
signal MULT_22:MULT_X;
signal MULT_23:MULT_X;
signal MULT_24:MULT_X;
signal MULT_25:MULT_X;
signal MULT_26:MULT_X;
signal MULT_27:MULT_X;
signal MULT_28:MULT_X;
signal MULT_29:MULT_X;
signal MULT_30:MULT_X;
signal MULT_31:MULT_X;
signal MULT_32:MULT_X;
signal MULT_33:MULT_X;
signal MULT_34:MULT_X;
signal MULT_35:MULT_X;
signal MULT_36:MULT_X;
signal MULT_37:MULT_X;
signal MULT_38:MULT_X;
signal MULT_39:MULT_X;
signal MULT_40:MULT_X;
signal MULT_41:MULT_X;
signal MULT_42:MULT_X;
signal MULT_43:MULT_X;
signal MULT_44:MULT_X;
signal MULT_45:MULT_X;
signal MULT_46:MULT_X;
signal MULT_47:MULT_X;
signal MULT_48:MULT_X;
signal MULT_49:MULT_X;
signal MULT_50:MULT_X;
signal MULT_51:MULT_X;
signal MULT_52:MULT_X;
signal MULT_53:MULT_X;
signal MULT_54:MULT_X;
signal MULT_55:MULT_X;
signal MULT_56:MULT_X;
signal MULT_57:MULT_X;
signal MULT_58:MULT_X;
signal MULT_59:MULT_X;
signal MULT_60:MULT_X;
signal MULT_61:MULT_X;
signal MULT_62:MULT_X;
signal MULT_63:MULT_X;
signal MULT_64:MULT_X;
signal MULT_65:MULT_X;
signal MULT_66:MULT_X;
signal MULT_67:MULT_X;
signal MULT_68:MULT_X;
signal MULT_69:MULT_X;
signal MULT_70:MULT_X;
signal MULT_71:MULT_X;
signal MULT_72:MULT_X;
signal MULT_73:MULT_X;
signal MULT_74:MULT_X;
signal MULT_75:MULT_X;
signal MULT_76:MULT_X;
signal MULT_77:MULT_X;
signal MULT_78:MULT_X;
signal MULT_79:MULT_X;
signal MULT_80:MULT_X;
signal MULT_81:MULT_X;
signal MULT_82:MULT_X;
signal MULT_83:MULT_X;
signal MULT_84:MULT_X;
signal DOUT_BUF_1_8	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_1		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_1		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_2_8	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_2		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_2		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_3_8	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_3		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_3		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_4_8	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_4		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_4		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_5_8	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_5		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_5		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_6_8	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_6		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_6		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_7_8	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_7		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_7		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_8_8	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_8		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_8		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_9_8	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_9		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_9		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_10_8	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_10		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_10		: signed(BIAS_SIZE-1   downto 0);


------------------------------------------------------ MULT SUMMATION DECLARATION-----------------------------------------------------------
signal SUM_PIXELS_1: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_2: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_3: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_4: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_5: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_6: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_7: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_8: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_9: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_10: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_11: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_12: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_13: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_14: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_15: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_16: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_17: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_18: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_19: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_20: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_21: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_22: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_23: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_24: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_25: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_26: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_27: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_28: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_29: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_30: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_31: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_32: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_33: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_34: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_35: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_36: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_37: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_38: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_39: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_40: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_41: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_42: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_43: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_44: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_45: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_46: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_47: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_48: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_49: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_50: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_51: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_52: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_53: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_54: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_55: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_56: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_57: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_58: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_59: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_60: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_61: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_62: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_63: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_64: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_65: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_66: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_67: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_68: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_69: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_70: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_71: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_72: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_73: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_74: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_75: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_76: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_77: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_78: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_79: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_80: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_81: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_82: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_83: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_84: signed(SUM_PEXILS-1 downto 0);
type    MULT_X_SUM_1	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_1- 1 downto 0);
signal  EN_SUM_MULT_1	: std_logic;
signal  MULTS_1_1:MULT_X_SUM_1;
signal  MULTS_1_2:MULT_X_SUM_1;
signal  MULTS_1_3:MULT_X_SUM_1;
signal  MULTS_1_4:MULT_X_SUM_1;
signal  MULTS_1_5:MULT_X_SUM_1;
signal  MULTS_1_6:MULT_X_SUM_1;
signal  MULTS_1_7:MULT_X_SUM_1;
signal  MULTS_1_8:MULT_X_SUM_1;
signal  MULTS_1_9:MULT_X_SUM_1;
signal  MULTS_1_10:MULT_X_SUM_1;
signal  MULTS_1_11:MULT_X_SUM_1;
signal  MULTS_1_12:MULT_X_SUM_1;
signal  MULTS_1_13:MULT_X_SUM_1;
signal  MULTS_1_14:MULT_X_SUM_1;
signal  MULTS_1_15:MULT_X_SUM_1;
signal  MULTS_1_16:MULT_X_SUM_1;
signal  MULTS_1_17:MULT_X_SUM_1;
signal  MULTS_1_18:MULT_X_SUM_1;
signal  MULTS_1_19:MULT_X_SUM_1;
signal  MULTS_1_20:MULT_X_SUM_1;
signal  MULTS_1_21:MULT_X_SUM_1;
signal  MULTS_1_22:MULT_X_SUM_1;
signal  MULTS_1_23:MULT_X_SUM_1;
signal  MULTS_1_24:MULT_X_SUM_1;
signal  MULTS_1_25:MULT_X_SUM_1;
signal  MULTS_1_26:MULT_X_SUM_1;
signal  MULTS_1_27:MULT_X_SUM_1;
signal  MULTS_1_28:MULT_X_SUM_1;
signal  MULTS_1_29:MULT_X_SUM_1;
signal  MULTS_1_30:MULT_X_SUM_1;
signal  MULTS_1_31:MULT_X_SUM_1;
signal  MULTS_1_32:MULT_X_SUM_1;
signal  MULTS_1_33:MULT_X_SUM_1;
signal  MULTS_1_34:MULT_X_SUM_1;
signal  MULTS_1_35:MULT_X_SUM_1;
signal  MULTS_1_36:MULT_X_SUM_1;
signal  MULTS_1_37:MULT_X_SUM_1;
signal  MULTS_1_38:MULT_X_SUM_1;
signal  MULTS_1_39:MULT_X_SUM_1;
signal  MULTS_1_40:MULT_X_SUM_1;
signal  MULTS_1_41:MULT_X_SUM_1;
signal  MULTS_1_42:MULT_X_SUM_1;
signal  MULTS_1_43:MULT_X_SUM_1;
signal  MULTS_1_44:MULT_X_SUM_1;
signal  MULTS_1_45:MULT_X_SUM_1;
signal  MULTS_1_46:MULT_X_SUM_1;
signal  MULTS_1_47:MULT_X_SUM_1;
signal  MULTS_1_48:MULT_X_SUM_1;
signal  MULTS_1_49:MULT_X_SUM_1;
signal  MULTS_1_50:MULT_X_SUM_1;
signal  MULTS_1_51:MULT_X_SUM_1;
signal  MULTS_1_52:MULT_X_SUM_1;
signal  MULTS_1_53:MULT_X_SUM_1;
signal  MULTS_1_54:MULT_X_SUM_1;
signal  MULTS_1_55:MULT_X_SUM_1;
signal  MULTS_1_56:MULT_X_SUM_1;
signal  MULTS_1_57:MULT_X_SUM_1;
signal  MULTS_1_58:MULT_X_SUM_1;
signal  MULTS_1_59:MULT_X_SUM_1;
signal  MULTS_1_60:MULT_X_SUM_1;
signal  MULTS_1_61:MULT_X_SUM_1;
signal  MULTS_1_62:MULT_X_SUM_1;
signal  MULTS_1_63:MULT_X_SUM_1;
signal  MULTS_1_64:MULT_X_SUM_1;
signal  MULTS_1_65:MULT_X_SUM_1;
signal  MULTS_1_66:MULT_X_SUM_1;
signal  MULTS_1_67:MULT_X_SUM_1;
signal  MULTS_1_68:MULT_X_SUM_1;
signal  MULTS_1_69:MULT_X_SUM_1;
signal  MULTS_1_70:MULT_X_SUM_1;
signal  MULTS_1_71:MULT_X_SUM_1;
signal  MULTS_1_72:MULT_X_SUM_1;
signal  MULTS_1_73:MULT_X_SUM_1;
signal  MULTS_1_74:MULT_X_SUM_1;
signal  MULTS_1_75:MULT_X_SUM_1;
signal  MULTS_1_76:MULT_X_SUM_1;
signal  MULTS_1_77:MULT_X_SUM_1;
signal  MULTS_1_78:MULT_X_SUM_1;
signal  MULTS_1_79:MULT_X_SUM_1;
signal  MULTS_1_80:MULT_X_SUM_1;
signal  MULTS_1_81:MULT_X_SUM_1;
signal  MULTS_1_82:MULT_X_SUM_1;
signal  MULTS_1_83:MULT_X_SUM_1;
signal  MULTS_1_84:MULT_X_SUM_1;
type    MULT_X_SUM_2	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_2- 1 downto 0);
signal  EN_SUM_MULT_2	: std_logic;
signal  MULTS_2_1:MULT_X_SUM_2;
signal  MULTS_2_2:MULT_X_SUM_2;
signal  MULTS_2_3:MULT_X_SUM_2;
signal  MULTS_2_4:MULT_X_SUM_2;
signal  MULTS_2_5:MULT_X_SUM_2;
signal  MULTS_2_6:MULT_X_SUM_2;
signal  MULTS_2_7:MULT_X_SUM_2;
signal  MULTS_2_8:MULT_X_SUM_2;
signal  MULTS_2_9:MULT_X_SUM_2;
signal  MULTS_2_10:MULT_X_SUM_2;
signal  MULTS_2_11:MULT_X_SUM_2;
signal  MULTS_2_12:MULT_X_SUM_2;
signal  MULTS_2_13:MULT_X_SUM_2;
signal  MULTS_2_14:MULT_X_SUM_2;
signal  MULTS_2_15:MULT_X_SUM_2;
signal  MULTS_2_16:MULT_X_SUM_2;
signal  MULTS_2_17:MULT_X_SUM_2;
signal  MULTS_2_18:MULT_X_SUM_2;
signal  MULTS_2_19:MULT_X_SUM_2;
signal  MULTS_2_20:MULT_X_SUM_2;
signal  MULTS_2_21:MULT_X_SUM_2;
signal  MULTS_2_22:MULT_X_SUM_2;
signal  MULTS_2_23:MULT_X_SUM_2;
signal  MULTS_2_24:MULT_X_SUM_2;
signal  MULTS_2_25:MULT_X_SUM_2;
signal  MULTS_2_26:MULT_X_SUM_2;
signal  MULTS_2_27:MULT_X_SUM_2;
signal  MULTS_2_28:MULT_X_SUM_2;
signal  MULTS_2_29:MULT_X_SUM_2;
signal  MULTS_2_30:MULT_X_SUM_2;
signal  MULTS_2_31:MULT_X_SUM_2;
signal  MULTS_2_32:MULT_X_SUM_2;
signal  MULTS_2_33:MULT_X_SUM_2;
signal  MULTS_2_34:MULT_X_SUM_2;
signal  MULTS_2_35:MULT_X_SUM_2;
signal  MULTS_2_36:MULT_X_SUM_2;
signal  MULTS_2_37:MULT_X_SUM_2;
signal  MULTS_2_38:MULT_X_SUM_2;
signal  MULTS_2_39:MULT_X_SUM_2;
signal  MULTS_2_40:MULT_X_SUM_2;
signal  MULTS_2_41:MULT_X_SUM_2;
signal  MULTS_2_42:MULT_X_SUM_2;
signal  MULTS_2_43:MULT_X_SUM_2;
signal  MULTS_2_44:MULT_X_SUM_2;
signal  MULTS_2_45:MULT_X_SUM_2;
signal  MULTS_2_46:MULT_X_SUM_2;
signal  MULTS_2_47:MULT_X_SUM_2;
signal  MULTS_2_48:MULT_X_SUM_2;
signal  MULTS_2_49:MULT_X_SUM_2;
signal  MULTS_2_50:MULT_X_SUM_2;
signal  MULTS_2_51:MULT_X_SUM_2;
signal  MULTS_2_52:MULT_X_SUM_2;
signal  MULTS_2_53:MULT_X_SUM_2;
signal  MULTS_2_54:MULT_X_SUM_2;
signal  MULTS_2_55:MULT_X_SUM_2;
signal  MULTS_2_56:MULT_X_SUM_2;
signal  MULTS_2_57:MULT_X_SUM_2;
signal  MULTS_2_58:MULT_X_SUM_2;
signal  MULTS_2_59:MULT_X_SUM_2;
signal  MULTS_2_60:MULT_X_SUM_2;
signal  MULTS_2_61:MULT_X_SUM_2;
signal  MULTS_2_62:MULT_X_SUM_2;
signal  MULTS_2_63:MULT_X_SUM_2;
signal  MULTS_2_64:MULT_X_SUM_2;
signal  MULTS_2_65:MULT_X_SUM_2;
signal  MULTS_2_66:MULT_X_SUM_2;
signal  MULTS_2_67:MULT_X_SUM_2;
signal  MULTS_2_68:MULT_X_SUM_2;
signal  MULTS_2_69:MULT_X_SUM_2;
signal  MULTS_2_70:MULT_X_SUM_2;
signal  MULTS_2_71:MULT_X_SUM_2;
signal  MULTS_2_72:MULT_X_SUM_2;
signal  MULTS_2_73:MULT_X_SUM_2;
signal  MULTS_2_74:MULT_X_SUM_2;
signal  MULTS_2_75:MULT_X_SUM_2;
signal  MULTS_2_76:MULT_X_SUM_2;
signal  MULTS_2_77:MULT_X_SUM_2;
signal  MULTS_2_78:MULT_X_SUM_2;
signal  MULTS_2_79:MULT_X_SUM_2;
signal  MULTS_2_80:MULT_X_SUM_2;
signal  MULTS_2_81:MULT_X_SUM_2;
signal  MULTS_2_82:MULT_X_SUM_2;
signal  MULTS_2_83:MULT_X_SUM_2;
signal  MULTS_2_84:MULT_X_SUM_2;
type    MULT_X_SUM_3	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_3- 1 downto 0);
signal  EN_SUM_MULT_3	: std_logic;
signal  MULTS_3_1:MULT_X_SUM_3;
signal  MULTS_3_2:MULT_X_SUM_3;
signal  MULTS_3_3:MULT_X_SUM_3;
signal  MULTS_3_4:MULT_X_SUM_3;
signal  MULTS_3_5:MULT_X_SUM_3;
signal  MULTS_3_6:MULT_X_SUM_3;
signal  MULTS_3_7:MULT_X_SUM_3;
signal  MULTS_3_8:MULT_X_SUM_3;
signal  MULTS_3_9:MULT_X_SUM_3;
signal  MULTS_3_10:MULT_X_SUM_3;
signal  MULTS_3_11:MULT_X_SUM_3;
signal  MULTS_3_12:MULT_X_SUM_3;
signal  MULTS_3_13:MULT_X_SUM_3;
signal  MULTS_3_14:MULT_X_SUM_3;
signal  MULTS_3_15:MULT_X_SUM_3;
signal  MULTS_3_16:MULT_X_SUM_3;
signal  MULTS_3_17:MULT_X_SUM_3;
signal  MULTS_3_18:MULT_X_SUM_3;
signal  MULTS_3_19:MULT_X_SUM_3;
signal  MULTS_3_20:MULT_X_SUM_3;
signal  MULTS_3_21:MULT_X_SUM_3;
signal  MULTS_3_22:MULT_X_SUM_3;
signal  MULTS_3_23:MULT_X_SUM_3;
signal  MULTS_3_24:MULT_X_SUM_3;
signal  MULTS_3_25:MULT_X_SUM_3;
signal  MULTS_3_26:MULT_X_SUM_3;
signal  MULTS_3_27:MULT_X_SUM_3;
signal  MULTS_3_28:MULT_X_SUM_3;
signal  MULTS_3_29:MULT_X_SUM_3;
signal  MULTS_3_30:MULT_X_SUM_3;
signal  MULTS_3_31:MULT_X_SUM_3;
signal  MULTS_3_32:MULT_X_SUM_3;
signal  MULTS_3_33:MULT_X_SUM_3;
signal  MULTS_3_34:MULT_X_SUM_3;
signal  MULTS_3_35:MULT_X_SUM_3;
signal  MULTS_3_36:MULT_X_SUM_3;
signal  MULTS_3_37:MULT_X_SUM_3;
signal  MULTS_3_38:MULT_X_SUM_3;
signal  MULTS_3_39:MULT_X_SUM_3;
signal  MULTS_3_40:MULT_X_SUM_3;
signal  MULTS_3_41:MULT_X_SUM_3;
signal  MULTS_3_42:MULT_X_SUM_3;
signal  MULTS_3_43:MULT_X_SUM_3;
signal  MULTS_3_44:MULT_X_SUM_3;
signal  MULTS_3_45:MULT_X_SUM_3;
signal  MULTS_3_46:MULT_X_SUM_3;
signal  MULTS_3_47:MULT_X_SUM_3;
signal  MULTS_3_48:MULT_X_SUM_3;
signal  MULTS_3_49:MULT_X_SUM_3;
signal  MULTS_3_50:MULT_X_SUM_3;
signal  MULTS_3_51:MULT_X_SUM_3;
signal  MULTS_3_52:MULT_X_SUM_3;
signal  MULTS_3_53:MULT_X_SUM_3;
signal  MULTS_3_54:MULT_X_SUM_3;
signal  MULTS_3_55:MULT_X_SUM_3;
signal  MULTS_3_56:MULT_X_SUM_3;
signal  MULTS_3_57:MULT_X_SUM_3;
signal  MULTS_3_58:MULT_X_SUM_3;
signal  MULTS_3_59:MULT_X_SUM_3;
signal  MULTS_3_60:MULT_X_SUM_3;
signal  MULTS_3_61:MULT_X_SUM_3;
signal  MULTS_3_62:MULT_X_SUM_3;
signal  MULTS_3_63:MULT_X_SUM_3;
signal  MULTS_3_64:MULT_X_SUM_3;
signal  MULTS_3_65:MULT_X_SUM_3;
signal  MULTS_3_66:MULT_X_SUM_3;
signal  MULTS_3_67:MULT_X_SUM_3;
signal  MULTS_3_68:MULT_X_SUM_3;
signal  MULTS_3_69:MULT_X_SUM_3;
signal  MULTS_3_70:MULT_X_SUM_3;
signal  MULTS_3_71:MULT_X_SUM_3;
signal  MULTS_3_72:MULT_X_SUM_3;
signal  MULTS_3_73:MULT_X_SUM_3;
signal  MULTS_3_74:MULT_X_SUM_3;
signal  MULTS_3_75:MULT_X_SUM_3;
signal  MULTS_3_76:MULT_X_SUM_3;
signal  MULTS_3_77:MULT_X_SUM_3;
signal  MULTS_3_78:MULT_X_SUM_3;
signal  MULTS_3_79:MULT_X_SUM_3;
signal  MULTS_3_80:MULT_X_SUM_3;
signal  MULTS_3_81:MULT_X_SUM_3;
signal  MULTS_3_82:MULT_X_SUM_3;
signal  MULTS_3_83:MULT_X_SUM_3;
signal  MULTS_3_84:MULT_X_SUM_3;
type    MULT_X_SUM_4	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_4- 1 downto 0);
signal  EN_SUM_MULT_4	: std_logic;
signal  MULTS_4_1:MULT_X_SUM_4;
signal  MULTS_4_2:MULT_X_SUM_4;
signal  MULTS_4_3:MULT_X_SUM_4;
signal  MULTS_4_4:MULT_X_SUM_4;
signal  MULTS_4_5:MULT_X_SUM_4;
signal  MULTS_4_6:MULT_X_SUM_4;
signal  MULTS_4_7:MULT_X_SUM_4;
signal  MULTS_4_8:MULT_X_SUM_4;
signal  MULTS_4_9:MULT_X_SUM_4;
signal  MULTS_4_10:MULT_X_SUM_4;
signal  MULTS_4_11:MULT_X_SUM_4;
signal  MULTS_4_12:MULT_X_SUM_4;
signal  MULTS_4_13:MULT_X_SUM_4;
signal  MULTS_4_14:MULT_X_SUM_4;
signal  MULTS_4_15:MULT_X_SUM_4;
signal  MULTS_4_16:MULT_X_SUM_4;
signal  MULTS_4_17:MULT_X_SUM_4;
signal  MULTS_4_18:MULT_X_SUM_4;
signal  MULTS_4_19:MULT_X_SUM_4;
signal  MULTS_4_20:MULT_X_SUM_4;
signal  MULTS_4_21:MULT_X_SUM_4;
signal  MULTS_4_22:MULT_X_SUM_4;
signal  MULTS_4_23:MULT_X_SUM_4;
signal  MULTS_4_24:MULT_X_SUM_4;
signal  MULTS_4_25:MULT_X_SUM_4;
signal  MULTS_4_26:MULT_X_SUM_4;
signal  MULTS_4_27:MULT_X_SUM_4;
signal  MULTS_4_28:MULT_X_SUM_4;
signal  MULTS_4_29:MULT_X_SUM_4;
signal  MULTS_4_30:MULT_X_SUM_4;
signal  MULTS_4_31:MULT_X_SUM_4;
signal  MULTS_4_32:MULT_X_SUM_4;
signal  MULTS_4_33:MULT_X_SUM_4;
signal  MULTS_4_34:MULT_X_SUM_4;
signal  MULTS_4_35:MULT_X_SUM_4;
signal  MULTS_4_36:MULT_X_SUM_4;
signal  MULTS_4_37:MULT_X_SUM_4;
signal  MULTS_4_38:MULT_X_SUM_4;
signal  MULTS_4_39:MULT_X_SUM_4;
signal  MULTS_4_40:MULT_X_SUM_4;
signal  MULTS_4_41:MULT_X_SUM_4;
signal  MULTS_4_42:MULT_X_SUM_4;
signal  MULTS_4_43:MULT_X_SUM_4;
signal  MULTS_4_44:MULT_X_SUM_4;
signal  MULTS_4_45:MULT_X_SUM_4;
signal  MULTS_4_46:MULT_X_SUM_4;
signal  MULTS_4_47:MULT_X_SUM_4;
signal  MULTS_4_48:MULT_X_SUM_4;
signal  MULTS_4_49:MULT_X_SUM_4;
signal  MULTS_4_50:MULT_X_SUM_4;
signal  MULTS_4_51:MULT_X_SUM_4;
signal  MULTS_4_52:MULT_X_SUM_4;
signal  MULTS_4_53:MULT_X_SUM_4;
signal  MULTS_4_54:MULT_X_SUM_4;
signal  MULTS_4_55:MULT_X_SUM_4;
signal  MULTS_4_56:MULT_X_SUM_4;
signal  MULTS_4_57:MULT_X_SUM_4;
signal  MULTS_4_58:MULT_X_SUM_4;
signal  MULTS_4_59:MULT_X_SUM_4;
signal  MULTS_4_60:MULT_X_SUM_4;
signal  MULTS_4_61:MULT_X_SUM_4;
signal  MULTS_4_62:MULT_X_SUM_4;
signal  MULTS_4_63:MULT_X_SUM_4;
signal  MULTS_4_64:MULT_X_SUM_4;
signal  MULTS_4_65:MULT_X_SUM_4;
signal  MULTS_4_66:MULT_X_SUM_4;
signal  MULTS_4_67:MULT_X_SUM_4;
signal  MULTS_4_68:MULT_X_SUM_4;
signal  MULTS_4_69:MULT_X_SUM_4;
signal  MULTS_4_70:MULT_X_SUM_4;
signal  MULTS_4_71:MULT_X_SUM_4;
signal  MULTS_4_72:MULT_X_SUM_4;
signal  MULTS_4_73:MULT_X_SUM_4;
signal  MULTS_4_74:MULT_X_SUM_4;
signal  MULTS_4_75:MULT_X_SUM_4;
signal  MULTS_4_76:MULT_X_SUM_4;
signal  MULTS_4_77:MULT_X_SUM_4;
signal  MULTS_4_78:MULT_X_SUM_4;
signal  MULTS_4_79:MULT_X_SUM_4;
signal  MULTS_4_80:MULT_X_SUM_4;
signal  MULTS_4_81:MULT_X_SUM_4;
signal  MULTS_4_82:MULT_X_SUM_4;
signal  MULTS_4_83:MULT_X_SUM_4;
signal  MULTS_4_84:MULT_X_SUM_4;
type    MULT_X_SUM_5	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_5- 1 downto 0);
signal  EN_SUM_MULT_5	: std_logic;
signal  MULTS_5_1:MULT_X_SUM_5;
signal  MULTS_5_2:MULT_X_SUM_5;
signal  MULTS_5_3:MULT_X_SUM_5;
signal  MULTS_5_4:MULT_X_SUM_5;
signal  MULTS_5_5:MULT_X_SUM_5;
signal  MULTS_5_6:MULT_X_SUM_5;
signal  MULTS_5_7:MULT_X_SUM_5;
signal  MULTS_5_8:MULT_X_SUM_5;
signal  MULTS_5_9:MULT_X_SUM_5;
signal  MULTS_5_10:MULT_X_SUM_5;
signal  MULTS_5_11:MULT_X_SUM_5;
signal  MULTS_5_12:MULT_X_SUM_5;
signal  MULTS_5_13:MULT_X_SUM_5;
signal  MULTS_5_14:MULT_X_SUM_5;
signal  MULTS_5_15:MULT_X_SUM_5;
signal  MULTS_5_16:MULT_X_SUM_5;
signal  MULTS_5_17:MULT_X_SUM_5;
signal  MULTS_5_18:MULT_X_SUM_5;
signal  MULTS_5_19:MULT_X_SUM_5;
signal  MULTS_5_20:MULT_X_SUM_5;
signal  MULTS_5_21:MULT_X_SUM_5;
signal  MULTS_5_22:MULT_X_SUM_5;
signal  MULTS_5_23:MULT_X_SUM_5;
signal  MULTS_5_24:MULT_X_SUM_5;
signal  MULTS_5_25:MULT_X_SUM_5;
signal  MULTS_5_26:MULT_X_SUM_5;
signal  MULTS_5_27:MULT_X_SUM_5;
signal  MULTS_5_28:MULT_X_SUM_5;
signal  MULTS_5_29:MULT_X_SUM_5;
signal  MULTS_5_30:MULT_X_SUM_5;
signal  MULTS_5_31:MULT_X_SUM_5;
signal  MULTS_5_32:MULT_X_SUM_5;
signal  MULTS_5_33:MULT_X_SUM_5;
signal  MULTS_5_34:MULT_X_SUM_5;
signal  MULTS_5_35:MULT_X_SUM_5;
signal  MULTS_5_36:MULT_X_SUM_5;
signal  MULTS_5_37:MULT_X_SUM_5;
signal  MULTS_5_38:MULT_X_SUM_5;
signal  MULTS_5_39:MULT_X_SUM_5;
signal  MULTS_5_40:MULT_X_SUM_5;
signal  MULTS_5_41:MULT_X_SUM_5;
signal  MULTS_5_42:MULT_X_SUM_5;
signal  MULTS_5_43:MULT_X_SUM_5;
signal  MULTS_5_44:MULT_X_SUM_5;
signal  MULTS_5_45:MULT_X_SUM_5;
signal  MULTS_5_46:MULT_X_SUM_5;
signal  MULTS_5_47:MULT_X_SUM_5;
signal  MULTS_5_48:MULT_X_SUM_5;
signal  MULTS_5_49:MULT_X_SUM_5;
signal  MULTS_5_50:MULT_X_SUM_5;
signal  MULTS_5_51:MULT_X_SUM_5;
signal  MULTS_5_52:MULT_X_SUM_5;
signal  MULTS_5_53:MULT_X_SUM_5;
signal  MULTS_5_54:MULT_X_SUM_5;
signal  MULTS_5_55:MULT_X_SUM_5;
signal  MULTS_5_56:MULT_X_SUM_5;
signal  MULTS_5_57:MULT_X_SUM_5;
signal  MULTS_5_58:MULT_X_SUM_5;
signal  MULTS_5_59:MULT_X_SUM_5;
signal  MULTS_5_60:MULT_X_SUM_5;
signal  MULTS_5_61:MULT_X_SUM_5;
signal  MULTS_5_62:MULT_X_SUM_5;
signal  MULTS_5_63:MULT_X_SUM_5;
signal  MULTS_5_64:MULT_X_SUM_5;
signal  MULTS_5_65:MULT_X_SUM_5;
signal  MULTS_5_66:MULT_X_SUM_5;
signal  MULTS_5_67:MULT_X_SUM_5;
signal  MULTS_5_68:MULT_X_SUM_5;
signal  MULTS_5_69:MULT_X_SUM_5;
signal  MULTS_5_70:MULT_X_SUM_5;
signal  MULTS_5_71:MULT_X_SUM_5;
signal  MULTS_5_72:MULT_X_SUM_5;
signal  MULTS_5_73:MULT_X_SUM_5;
signal  MULTS_5_74:MULT_X_SUM_5;
signal  MULTS_5_75:MULT_X_SUM_5;
signal  MULTS_5_76:MULT_X_SUM_5;
signal  MULTS_5_77:MULT_X_SUM_5;
signal  MULTS_5_78:MULT_X_SUM_5;
signal  MULTS_5_79:MULT_X_SUM_5;
signal  MULTS_5_80:MULT_X_SUM_5;
signal  MULTS_5_81:MULT_X_SUM_5;
signal  MULTS_5_82:MULT_X_SUM_5;
signal  MULTS_5_83:MULT_X_SUM_5;
signal  MULTS_5_84:MULT_X_SUM_5;
type    MULT_X_SUM_6	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_6- 1 downto 0);
signal  EN_SUM_MULT_6	: std_logic;
signal  MULTS_6_1:MULT_X_SUM_6;
signal  MULTS_6_2:MULT_X_SUM_6;
signal  MULTS_6_3:MULT_X_SUM_6;
signal  MULTS_6_4:MULT_X_SUM_6;
signal  MULTS_6_5:MULT_X_SUM_6;
signal  MULTS_6_6:MULT_X_SUM_6;
signal  MULTS_6_7:MULT_X_SUM_6;
signal  MULTS_6_8:MULT_X_SUM_6;
signal  MULTS_6_9:MULT_X_SUM_6;
signal  MULTS_6_10:MULT_X_SUM_6;
signal  MULTS_6_11:MULT_X_SUM_6;
signal  MULTS_6_12:MULT_X_SUM_6;
signal  MULTS_6_13:MULT_X_SUM_6;
signal  MULTS_6_14:MULT_X_SUM_6;
signal  MULTS_6_15:MULT_X_SUM_6;
signal  MULTS_6_16:MULT_X_SUM_6;
signal  MULTS_6_17:MULT_X_SUM_6;
signal  MULTS_6_18:MULT_X_SUM_6;
signal  MULTS_6_19:MULT_X_SUM_6;
signal  MULTS_6_20:MULT_X_SUM_6;
signal  MULTS_6_21:MULT_X_SUM_6;
signal  MULTS_6_22:MULT_X_SUM_6;
signal  MULTS_6_23:MULT_X_SUM_6;
signal  MULTS_6_24:MULT_X_SUM_6;
signal  MULTS_6_25:MULT_X_SUM_6;
signal  MULTS_6_26:MULT_X_SUM_6;
signal  MULTS_6_27:MULT_X_SUM_6;
signal  MULTS_6_28:MULT_X_SUM_6;
signal  MULTS_6_29:MULT_X_SUM_6;
signal  MULTS_6_30:MULT_X_SUM_6;
signal  MULTS_6_31:MULT_X_SUM_6;
signal  MULTS_6_32:MULT_X_SUM_6;
signal  MULTS_6_33:MULT_X_SUM_6;
signal  MULTS_6_34:MULT_X_SUM_6;
signal  MULTS_6_35:MULT_X_SUM_6;
signal  MULTS_6_36:MULT_X_SUM_6;
signal  MULTS_6_37:MULT_X_SUM_6;
signal  MULTS_6_38:MULT_X_SUM_6;
signal  MULTS_6_39:MULT_X_SUM_6;
signal  MULTS_6_40:MULT_X_SUM_6;
signal  MULTS_6_41:MULT_X_SUM_6;
signal  MULTS_6_42:MULT_X_SUM_6;
signal  MULTS_6_43:MULT_X_SUM_6;
signal  MULTS_6_44:MULT_X_SUM_6;
signal  MULTS_6_45:MULT_X_SUM_6;
signal  MULTS_6_46:MULT_X_SUM_6;
signal  MULTS_6_47:MULT_X_SUM_6;
signal  MULTS_6_48:MULT_X_SUM_6;
signal  MULTS_6_49:MULT_X_SUM_6;
signal  MULTS_6_50:MULT_X_SUM_6;
signal  MULTS_6_51:MULT_X_SUM_6;
signal  MULTS_6_52:MULT_X_SUM_6;
signal  MULTS_6_53:MULT_X_SUM_6;
signal  MULTS_6_54:MULT_X_SUM_6;
signal  MULTS_6_55:MULT_X_SUM_6;
signal  MULTS_6_56:MULT_X_SUM_6;
signal  MULTS_6_57:MULT_X_SUM_6;
signal  MULTS_6_58:MULT_X_SUM_6;
signal  MULTS_6_59:MULT_X_SUM_6;
signal  MULTS_6_60:MULT_X_SUM_6;
signal  MULTS_6_61:MULT_X_SUM_6;
signal  MULTS_6_62:MULT_X_SUM_6;
signal  MULTS_6_63:MULT_X_SUM_6;
signal  MULTS_6_64:MULT_X_SUM_6;
signal  MULTS_6_65:MULT_X_SUM_6;
signal  MULTS_6_66:MULT_X_SUM_6;
signal  MULTS_6_67:MULT_X_SUM_6;
signal  MULTS_6_68:MULT_X_SUM_6;
signal  MULTS_6_69:MULT_X_SUM_6;
signal  MULTS_6_70:MULT_X_SUM_6;
signal  MULTS_6_71:MULT_X_SUM_6;
signal  MULTS_6_72:MULT_X_SUM_6;
signal  MULTS_6_73:MULT_X_SUM_6;
signal  MULTS_6_74:MULT_X_SUM_6;
signal  MULTS_6_75:MULT_X_SUM_6;
signal  MULTS_6_76:MULT_X_SUM_6;
signal  MULTS_6_77:MULT_X_SUM_6;
signal  MULTS_6_78:MULT_X_SUM_6;
signal  MULTS_6_79:MULT_X_SUM_6;
signal  MULTS_6_80:MULT_X_SUM_6;
signal  MULTS_6_81:MULT_X_SUM_6;
signal  MULTS_6_82:MULT_X_SUM_6;
signal  MULTS_6_83:MULT_X_SUM_6;
signal  MULTS_6_84:MULT_X_SUM_6;
type    MULT_X_SUM_7	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_7- 1 downto 0);
signal  EN_SUM_MULT_7	: std_logic;
signal  MULTS_7_1:MULT_X_SUM_7;
signal  MULTS_7_2:MULT_X_SUM_7;
signal  MULTS_7_3:MULT_X_SUM_7;
signal  MULTS_7_4:MULT_X_SUM_7;
signal  MULTS_7_5:MULT_X_SUM_7;
signal  MULTS_7_6:MULT_X_SUM_7;
signal  MULTS_7_7:MULT_X_SUM_7;
signal  MULTS_7_8:MULT_X_SUM_7;
signal  MULTS_7_9:MULT_X_SUM_7;
signal  MULTS_7_10:MULT_X_SUM_7;
signal  MULTS_7_11:MULT_X_SUM_7;
signal  MULTS_7_12:MULT_X_SUM_7;
signal  MULTS_7_13:MULT_X_SUM_7;
signal  MULTS_7_14:MULT_X_SUM_7;
signal  MULTS_7_15:MULT_X_SUM_7;
signal  MULTS_7_16:MULT_X_SUM_7;
signal  MULTS_7_17:MULT_X_SUM_7;
signal  MULTS_7_18:MULT_X_SUM_7;
signal  MULTS_7_19:MULT_X_SUM_7;
signal  MULTS_7_20:MULT_X_SUM_7;
signal  MULTS_7_21:MULT_X_SUM_7;
signal  MULTS_7_22:MULT_X_SUM_7;
signal  MULTS_7_23:MULT_X_SUM_7;
signal  MULTS_7_24:MULT_X_SUM_7;
signal  MULTS_7_25:MULT_X_SUM_7;
signal  MULTS_7_26:MULT_X_SUM_7;
signal  MULTS_7_27:MULT_X_SUM_7;
signal  MULTS_7_28:MULT_X_SUM_7;
signal  MULTS_7_29:MULT_X_SUM_7;
signal  MULTS_7_30:MULT_X_SUM_7;
signal  MULTS_7_31:MULT_X_SUM_7;
signal  MULTS_7_32:MULT_X_SUM_7;
signal  MULTS_7_33:MULT_X_SUM_7;
signal  MULTS_7_34:MULT_X_SUM_7;
signal  MULTS_7_35:MULT_X_SUM_7;
signal  MULTS_7_36:MULT_X_SUM_7;
signal  MULTS_7_37:MULT_X_SUM_7;
signal  MULTS_7_38:MULT_X_SUM_7;
signal  MULTS_7_39:MULT_X_SUM_7;
signal  MULTS_7_40:MULT_X_SUM_7;
signal  MULTS_7_41:MULT_X_SUM_7;
signal  MULTS_7_42:MULT_X_SUM_7;
signal  MULTS_7_43:MULT_X_SUM_7;
signal  MULTS_7_44:MULT_X_SUM_7;
signal  MULTS_7_45:MULT_X_SUM_7;
signal  MULTS_7_46:MULT_X_SUM_7;
signal  MULTS_7_47:MULT_X_SUM_7;
signal  MULTS_7_48:MULT_X_SUM_7;
signal  MULTS_7_49:MULT_X_SUM_7;
signal  MULTS_7_50:MULT_X_SUM_7;
signal  MULTS_7_51:MULT_X_SUM_7;
signal  MULTS_7_52:MULT_X_SUM_7;
signal  MULTS_7_53:MULT_X_SUM_7;
signal  MULTS_7_54:MULT_X_SUM_7;
signal  MULTS_7_55:MULT_X_SUM_7;
signal  MULTS_7_56:MULT_X_SUM_7;
signal  MULTS_7_57:MULT_X_SUM_7;
signal  MULTS_7_58:MULT_X_SUM_7;
signal  MULTS_7_59:MULT_X_SUM_7;
signal  MULTS_7_60:MULT_X_SUM_7;
signal  MULTS_7_61:MULT_X_SUM_7;
signal  MULTS_7_62:MULT_X_SUM_7;
signal  MULTS_7_63:MULT_X_SUM_7;
signal  MULTS_7_64:MULT_X_SUM_7;
signal  MULTS_7_65:MULT_X_SUM_7;
signal  MULTS_7_66:MULT_X_SUM_7;
signal  MULTS_7_67:MULT_X_SUM_7;
signal  MULTS_7_68:MULT_X_SUM_7;
signal  MULTS_7_69:MULT_X_SUM_7;
signal  MULTS_7_70:MULT_X_SUM_7;
signal  MULTS_7_71:MULT_X_SUM_7;
signal  MULTS_7_72:MULT_X_SUM_7;
signal  MULTS_7_73:MULT_X_SUM_7;
signal  MULTS_7_74:MULT_X_SUM_7;
signal  MULTS_7_75:MULT_X_SUM_7;
signal  MULTS_7_76:MULT_X_SUM_7;
signal  MULTS_7_77:MULT_X_SUM_7;
signal  MULTS_7_78:MULT_X_SUM_7;
signal  MULTS_7_79:MULT_X_SUM_7;
signal  MULTS_7_80:MULT_X_SUM_7;
signal  MULTS_7_81:MULT_X_SUM_7;
signal  MULTS_7_82:MULT_X_SUM_7;
signal  MULTS_7_83:MULT_X_SUM_7;
signal  MULTS_7_84:MULT_X_SUM_7;



--------------------------------------------- FILTER HARDCODED CONSTANTS -WEIGHTS START--------------------------------

constant FMAP_1_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";

constant BIAS_VAL_1: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_2: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_3: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_4: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_5: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_6: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_7: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_8: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_9: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_10: signed (BIASES_SIZE-1 downto 0):="01";


BEGIN
-------------------------------------------------------- ARCHITECTURE BEGIN--------------------------------------------------------

LAYER_8: process(CLK)


begin
------------------------------------------------ RESET AND PROCESS TOP START ------------------------------------------------------
if rising_edge(CLK) then
  if RST = '1' then
	-------------------FIXED SIGNALS RESET------------------------
    PIXEL_COUNT<=0;VALID_NXTLYR_PIX<=0;OUT_PIXEL_COUNT<=0;
    EN_NXT_LYR_8<='0';FRST_TIM_EN_8<='0';INTERNAL_RST<='0';
    Enable_MULT<='0';Enable_ADDER<='0';Enable_ReLU<='0';Enable_BIAS<='0';
    PADDING_count<=0;ROW_COUNT<=0;SIG_STRIDE<=STRIDE;COUNT_PIX<=0;

-------------------DYNAMIC SIGNALS RESET------------------------
    DOUT_BUF_1_8<=(others => '0');BIAS_1<=(others => '0');ReLU_1<=(others => '0');
    DOUT_BUF_2_8<=(others => '0');BIAS_2<=(others => '0');ReLU_2<=(others => '0');
    DOUT_BUF_3_8<=(others => '0');BIAS_3<=(others => '0');ReLU_3<=(others => '0');
    DOUT_BUF_4_8<=(others => '0');BIAS_4<=(others => '0');ReLU_4<=(others => '0');
    DOUT_BUF_5_8<=(others => '0');BIAS_5<=(others => '0');ReLU_5<=(others => '0');
    DOUT_BUF_6_8<=(others => '0');BIAS_6<=(others => '0');ReLU_6<=(others => '0');
    DOUT_BUF_7_8<=(others => '0');BIAS_7<=(others => '0');ReLU_7<=(others => '0');
    DOUT_BUF_8_8<=(others => '0');BIAS_8<=(others => '0');ReLU_8<=(others => '0');
    DOUT_BUF_9_8<=(others => '0');BIAS_9<=(others => '0');ReLU_9<=(others => '0');
    DOUT_BUF_10_8<=(others => '0');BIAS_10<=(others => '0');ReLU_10<=(others => '0');

    SUM_PIXELS_1<=(others=>'0');MULT_1<=((others=> (others=>'0')));
    SUM_PIXELS_2<=(others=>'0');MULT_2<=((others=> (others=>'0')));
    SUM_PIXELS_3<=(others=>'0');MULT_3<=((others=> (others=>'0')));
    SUM_PIXELS_4<=(others=>'0');MULT_4<=((others=> (others=>'0')));
    SUM_PIXELS_5<=(others=>'0');MULT_5<=((others=> (others=>'0')));
    SUM_PIXELS_6<=(others=>'0');MULT_6<=((others=> (others=>'0')));
    SUM_PIXELS_7<=(others=>'0');MULT_7<=((others=> (others=>'0')));
    SUM_PIXELS_8<=(others=>'0');MULT_8<=((others=> (others=>'0')));
    SUM_PIXELS_9<=(others=>'0');MULT_9<=((others=> (others=>'0')));
    SUM_PIXELS_10<=(others=>'0');MULT_10<=((others=> (others=>'0')));
    SUM_PIXELS_11<=(others=>'0');MULT_11<=((others=> (others=>'0')));
    SUM_PIXELS_12<=(others=>'0');MULT_12<=((others=> (others=>'0')));
    SUM_PIXELS_13<=(others=>'0');MULT_13<=((others=> (others=>'0')));
    SUM_PIXELS_14<=(others=>'0');MULT_14<=((others=> (others=>'0')));
    SUM_PIXELS_15<=(others=>'0');MULT_15<=((others=> (others=>'0')));
    SUM_PIXELS_16<=(others=>'0');MULT_16<=((others=> (others=>'0')));
    SUM_PIXELS_17<=(others=>'0');MULT_17<=((others=> (others=>'0')));
    SUM_PIXELS_18<=(others=>'0');MULT_18<=((others=> (others=>'0')));
    SUM_PIXELS_19<=(others=>'0');MULT_19<=((others=> (others=>'0')));
    SUM_PIXELS_20<=(others=>'0');MULT_20<=((others=> (others=>'0')));
    SUM_PIXELS_21<=(others=>'0');MULT_21<=((others=> (others=>'0')));
    SUM_PIXELS_22<=(others=>'0');MULT_22<=((others=> (others=>'0')));
    SUM_PIXELS_23<=(others=>'0');MULT_23<=((others=> (others=>'0')));
    SUM_PIXELS_24<=(others=>'0');MULT_24<=((others=> (others=>'0')));
    SUM_PIXELS_25<=(others=>'0');MULT_25<=((others=> (others=>'0')));
    SUM_PIXELS_26<=(others=>'0');MULT_26<=((others=> (others=>'0')));
    SUM_PIXELS_27<=(others=>'0');MULT_27<=((others=> (others=>'0')));
    SUM_PIXELS_28<=(others=>'0');MULT_28<=((others=> (others=>'0')));
    SUM_PIXELS_29<=(others=>'0');MULT_29<=((others=> (others=>'0')));
    SUM_PIXELS_30<=(others=>'0');MULT_30<=((others=> (others=>'0')));
    SUM_PIXELS_31<=(others=>'0');MULT_31<=((others=> (others=>'0')));
    SUM_PIXELS_32<=(others=>'0');MULT_32<=((others=> (others=>'0')));
    SUM_PIXELS_33<=(others=>'0');MULT_33<=((others=> (others=>'0')));
    SUM_PIXELS_34<=(others=>'0');MULT_34<=((others=> (others=>'0')));
    SUM_PIXELS_35<=(others=>'0');MULT_35<=((others=> (others=>'0')));
    SUM_PIXELS_36<=(others=>'0');MULT_36<=((others=> (others=>'0')));
    SUM_PIXELS_37<=(others=>'0');MULT_37<=((others=> (others=>'0')));
    SUM_PIXELS_38<=(others=>'0');MULT_38<=((others=> (others=>'0')));
    SUM_PIXELS_39<=(others=>'0');MULT_39<=((others=> (others=>'0')));
    SUM_PIXELS_40<=(others=>'0');MULT_40<=((others=> (others=>'0')));
    SUM_PIXELS_41<=(others=>'0');MULT_41<=((others=> (others=>'0')));
    SUM_PIXELS_42<=(others=>'0');MULT_42<=((others=> (others=>'0')));
    SUM_PIXELS_43<=(others=>'0');MULT_43<=((others=> (others=>'0')));
    SUM_PIXELS_44<=(others=>'0');MULT_44<=((others=> (others=>'0')));
    SUM_PIXELS_45<=(others=>'0');MULT_45<=((others=> (others=>'0')));
    SUM_PIXELS_46<=(others=>'0');MULT_46<=((others=> (others=>'0')));
    SUM_PIXELS_47<=(others=>'0');MULT_47<=((others=> (others=>'0')));
    SUM_PIXELS_48<=(others=>'0');MULT_48<=((others=> (others=>'0')));
    SUM_PIXELS_49<=(others=>'0');MULT_49<=((others=> (others=>'0')));
    SUM_PIXELS_50<=(others=>'0');MULT_50<=((others=> (others=>'0')));
    SUM_PIXELS_51<=(others=>'0');MULT_51<=((others=> (others=>'0')));
    SUM_PIXELS_52<=(others=>'0');MULT_52<=((others=> (others=>'0')));
    SUM_PIXELS_53<=(others=>'0');MULT_53<=((others=> (others=>'0')));
    SUM_PIXELS_54<=(others=>'0');MULT_54<=((others=> (others=>'0')));
    SUM_PIXELS_55<=(others=>'0');MULT_55<=((others=> (others=>'0')));
    SUM_PIXELS_56<=(others=>'0');MULT_56<=((others=> (others=>'0')));
    SUM_PIXELS_57<=(others=>'0');MULT_57<=((others=> (others=>'0')));
    SUM_PIXELS_58<=(others=>'0');MULT_58<=((others=> (others=>'0')));
    SUM_PIXELS_59<=(others=>'0');MULT_59<=((others=> (others=>'0')));
    SUM_PIXELS_60<=(others=>'0');MULT_60<=((others=> (others=>'0')));
    SUM_PIXELS_61<=(others=>'0');MULT_61<=((others=> (others=>'0')));
    SUM_PIXELS_62<=(others=>'0');MULT_62<=((others=> (others=>'0')));
    SUM_PIXELS_63<=(others=>'0');MULT_63<=((others=> (others=>'0')));
    SUM_PIXELS_64<=(others=>'0');MULT_64<=((others=> (others=>'0')));
    SUM_PIXELS_65<=(others=>'0');MULT_65<=((others=> (others=>'0')));
    SUM_PIXELS_66<=(others=>'0');MULT_66<=((others=> (others=>'0')));
    SUM_PIXELS_67<=(others=>'0');MULT_67<=((others=> (others=>'0')));
    SUM_PIXELS_68<=(others=>'0');MULT_68<=((others=> (others=>'0')));
    SUM_PIXELS_69<=(others=>'0');MULT_69<=((others=> (others=>'0')));
    SUM_PIXELS_70<=(others=>'0');MULT_70<=((others=> (others=>'0')));
    SUM_PIXELS_71<=(others=>'0');MULT_71<=((others=> (others=>'0')));
    SUM_PIXELS_72<=(others=>'0');MULT_72<=((others=> (others=>'0')));
    SUM_PIXELS_73<=(others=>'0');MULT_73<=((others=> (others=>'0')));
    SUM_PIXELS_74<=(others=>'0');MULT_74<=((others=> (others=>'0')));
    SUM_PIXELS_75<=(others=>'0');MULT_75<=((others=> (others=>'0')));
    SUM_PIXELS_76<=(others=>'0');MULT_76<=((others=> (others=>'0')));
    SUM_PIXELS_77<=(others=>'0');MULT_77<=((others=> (others=>'0')));
    SUM_PIXELS_78<=(others=>'0');MULT_78<=((others=> (others=>'0')));
    SUM_PIXELS_79<=(others=>'0');MULT_79<=((others=> (others=>'0')));
    SUM_PIXELS_80<=(others=>'0');MULT_80<=((others=> (others=>'0')));
    SUM_PIXELS_81<=(others=>'0');MULT_81<=((others=> (others=>'0')));
    SUM_PIXELS_82<=(others=>'0');MULT_82<=((others=> (others=>'0')));
    SUM_PIXELS_83<=(others=>'0');MULT_83<=((others=> (others=>'0')));
    SUM_PIXELS_84<=(others=>'0');MULT_84<=((others=> (others=>'0')));

    EN_SUM_MULT_1<='0';
    MULTS_1_1<=((others=> (others=>'0')));
    MULTS_1_2<=((others=> (others=>'0')));
    MULTS_1_3<=((others=> (others=>'0')));
    MULTS_1_4<=((others=> (others=>'0')));
    MULTS_1_5<=((others=> (others=>'0')));
    MULTS_1_6<=((others=> (others=>'0')));
    MULTS_1_7<=((others=> (others=>'0')));
    MULTS_1_8<=((others=> (others=>'0')));
    MULTS_1_9<=((others=> (others=>'0')));
    MULTS_1_10<=((others=> (others=>'0')));
    MULTS_1_11<=((others=> (others=>'0')));
    MULTS_1_12<=((others=> (others=>'0')));
    MULTS_1_13<=((others=> (others=>'0')));
    MULTS_1_14<=((others=> (others=>'0')));
    MULTS_1_15<=((others=> (others=>'0')));
    MULTS_1_16<=((others=> (others=>'0')));
    MULTS_1_17<=((others=> (others=>'0')));
    MULTS_1_18<=((others=> (others=>'0')));
    MULTS_1_19<=((others=> (others=>'0')));
    MULTS_1_20<=((others=> (others=>'0')));
    MULTS_1_21<=((others=> (others=>'0')));
    MULTS_1_22<=((others=> (others=>'0')));
    MULTS_1_23<=((others=> (others=>'0')));
    MULTS_1_24<=((others=> (others=>'0')));
    MULTS_1_25<=((others=> (others=>'0')));
    MULTS_1_26<=((others=> (others=>'0')));
    MULTS_1_27<=((others=> (others=>'0')));
    MULTS_1_28<=((others=> (others=>'0')));
    MULTS_1_29<=((others=> (others=>'0')));
    MULTS_1_30<=((others=> (others=>'0')));
    MULTS_1_31<=((others=> (others=>'0')));
    MULTS_1_32<=((others=> (others=>'0')));
    MULTS_1_33<=((others=> (others=>'0')));
    MULTS_1_34<=((others=> (others=>'0')));
    MULTS_1_35<=((others=> (others=>'0')));
    MULTS_1_36<=((others=> (others=>'0')));
    MULTS_1_37<=((others=> (others=>'0')));
    MULTS_1_38<=((others=> (others=>'0')));
    MULTS_1_39<=((others=> (others=>'0')));
    MULTS_1_40<=((others=> (others=>'0')));
    MULTS_1_41<=((others=> (others=>'0')));
    MULTS_1_42<=((others=> (others=>'0')));
    MULTS_1_43<=((others=> (others=>'0')));
    MULTS_1_44<=((others=> (others=>'0')));
    MULTS_1_45<=((others=> (others=>'0')));
    MULTS_1_46<=((others=> (others=>'0')));
    MULTS_1_47<=((others=> (others=>'0')));
    MULTS_1_48<=((others=> (others=>'0')));
    MULTS_1_49<=((others=> (others=>'0')));
    MULTS_1_50<=((others=> (others=>'0')));
    MULTS_1_51<=((others=> (others=>'0')));
    MULTS_1_52<=((others=> (others=>'0')));
    MULTS_1_53<=((others=> (others=>'0')));
    MULTS_1_54<=((others=> (others=>'0')));
    MULTS_1_55<=((others=> (others=>'0')));
    MULTS_1_56<=((others=> (others=>'0')));
    MULTS_1_57<=((others=> (others=>'0')));
    MULTS_1_58<=((others=> (others=>'0')));
    MULTS_1_59<=((others=> (others=>'0')));
    MULTS_1_60<=((others=> (others=>'0')));
    MULTS_1_61<=((others=> (others=>'0')));
    MULTS_1_62<=((others=> (others=>'0')));
    MULTS_1_63<=((others=> (others=>'0')));
    MULTS_1_64<=((others=> (others=>'0')));
    MULTS_1_65<=((others=> (others=>'0')));
    MULTS_1_66<=((others=> (others=>'0')));
    MULTS_1_67<=((others=> (others=>'0')));
    MULTS_1_68<=((others=> (others=>'0')));
    MULTS_1_69<=((others=> (others=>'0')));
    MULTS_1_70<=((others=> (others=>'0')));
    MULTS_1_71<=((others=> (others=>'0')));
    MULTS_1_72<=((others=> (others=>'0')));
    MULTS_1_73<=((others=> (others=>'0')));
    MULTS_1_74<=((others=> (others=>'0')));
    MULTS_1_75<=((others=> (others=>'0')));
    MULTS_1_76<=((others=> (others=>'0')));
    MULTS_1_77<=((others=> (others=>'0')));
    MULTS_1_78<=((others=> (others=>'0')));
    MULTS_1_79<=((others=> (others=>'0')));
    MULTS_1_80<=((others=> (others=>'0')));
    MULTS_1_81<=((others=> (others=>'0')));
    MULTS_1_82<=((others=> (others=>'0')));
    MULTS_1_83<=((others=> (others=>'0')));
    MULTS_1_84<=((others=> (others=>'0')));
    EN_SUM_MULT_2<='0';
    MULTS_2_1<=((others=> (others=>'0')));
    MULTS_2_2<=((others=> (others=>'0')));
    MULTS_2_3<=((others=> (others=>'0')));
    MULTS_2_4<=((others=> (others=>'0')));
    MULTS_2_5<=((others=> (others=>'0')));
    MULTS_2_6<=((others=> (others=>'0')));
    MULTS_2_7<=((others=> (others=>'0')));
    MULTS_2_8<=((others=> (others=>'0')));
    MULTS_2_9<=((others=> (others=>'0')));
    MULTS_2_10<=((others=> (others=>'0')));
    MULTS_2_11<=((others=> (others=>'0')));
    MULTS_2_12<=((others=> (others=>'0')));
    MULTS_2_13<=((others=> (others=>'0')));
    MULTS_2_14<=((others=> (others=>'0')));
    MULTS_2_15<=((others=> (others=>'0')));
    MULTS_2_16<=((others=> (others=>'0')));
    MULTS_2_17<=((others=> (others=>'0')));
    MULTS_2_18<=((others=> (others=>'0')));
    MULTS_2_19<=((others=> (others=>'0')));
    MULTS_2_20<=((others=> (others=>'0')));
    MULTS_2_21<=((others=> (others=>'0')));
    MULTS_2_22<=((others=> (others=>'0')));
    MULTS_2_23<=((others=> (others=>'0')));
    MULTS_2_24<=((others=> (others=>'0')));
    MULTS_2_25<=((others=> (others=>'0')));
    MULTS_2_26<=((others=> (others=>'0')));
    MULTS_2_27<=((others=> (others=>'0')));
    MULTS_2_28<=((others=> (others=>'0')));
    MULTS_2_29<=((others=> (others=>'0')));
    MULTS_2_30<=((others=> (others=>'0')));
    MULTS_2_31<=((others=> (others=>'0')));
    MULTS_2_32<=((others=> (others=>'0')));
    MULTS_2_33<=((others=> (others=>'0')));
    MULTS_2_34<=((others=> (others=>'0')));
    MULTS_2_35<=((others=> (others=>'0')));
    MULTS_2_36<=((others=> (others=>'0')));
    MULTS_2_37<=((others=> (others=>'0')));
    MULTS_2_38<=((others=> (others=>'0')));
    MULTS_2_39<=((others=> (others=>'0')));
    MULTS_2_40<=((others=> (others=>'0')));
    MULTS_2_41<=((others=> (others=>'0')));
    MULTS_2_42<=((others=> (others=>'0')));
    MULTS_2_43<=((others=> (others=>'0')));
    MULTS_2_44<=((others=> (others=>'0')));
    MULTS_2_45<=((others=> (others=>'0')));
    MULTS_2_46<=((others=> (others=>'0')));
    MULTS_2_47<=((others=> (others=>'0')));
    MULTS_2_48<=((others=> (others=>'0')));
    MULTS_2_49<=((others=> (others=>'0')));
    MULTS_2_50<=((others=> (others=>'0')));
    MULTS_2_51<=((others=> (others=>'0')));
    MULTS_2_52<=((others=> (others=>'0')));
    MULTS_2_53<=((others=> (others=>'0')));
    MULTS_2_54<=((others=> (others=>'0')));
    MULTS_2_55<=((others=> (others=>'0')));
    MULTS_2_56<=((others=> (others=>'0')));
    MULTS_2_57<=((others=> (others=>'0')));
    MULTS_2_58<=((others=> (others=>'0')));
    MULTS_2_59<=((others=> (others=>'0')));
    MULTS_2_60<=((others=> (others=>'0')));
    MULTS_2_61<=((others=> (others=>'0')));
    MULTS_2_62<=((others=> (others=>'0')));
    MULTS_2_63<=((others=> (others=>'0')));
    MULTS_2_64<=((others=> (others=>'0')));
    MULTS_2_65<=((others=> (others=>'0')));
    MULTS_2_66<=((others=> (others=>'0')));
    MULTS_2_67<=((others=> (others=>'0')));
    MULTS_2_68<=((others=> (others=>'0')));
    MULTS_2_69<=((others=> (others=>'0')));
    MULTS_2_70<=((others=> (others=>'0')));
    MULTS_2_71<=((others=> (others=>'0')));
    MULTS_2_72<=((others=> (others=>'0')));
    MULTS_2_73<=((others=> (others=>'0')));
    MULTS_2_74<=((others=> (others=>'0')));
    MULTS_2_75<=((others=> (others=>'0')));
    MULTS_2_76<=((others=> (others=>'0')));
    MULTS_2_77<=((others=> (others=>'0')));
    MULTS_2_78<=((others=> (others=>'0')));
    MULTS_2_79<=((others=> (others=>'0')));
    MULTS_2_80<=((others=> (others=>'0')));
    MULTS_2_81<=((others=> (others=>'0')));
    MULTS_2_82<=((others=> (others=>'0')));
    MULTS_2_83<=((others=> (others=>'0')));
    MULTS_2_84<=((others=> (others=>'0')));
    EN_SUM_MULT_3<='0';
    MULTS_3_1<=((others=> (others=>'0')));
    MULTS_3_2<=((others=> (others=>'0')));
    MULTS_3_3<=((others=> (others=>'0')));
    MULTS_3_4<=((others=> (others=>'0')));
    MULTS_3_5<=((others=> (others=>'0')));
    MULTS_3_6<=((others=> (others=>'0')));
    MULTS_3_7<=((others=> (others=>'0')));
    MULTS_3_8<=((others=> (others=>'0')));
    MULTS_3_9<=((others=> (others=>'0')));
    MULTS_3_10<=((others=> (others=>'0')));
    MULTS_3_11<=((others=> (others=>'0')));
    MULTS_3_12<=((others=> (others=>'0')));
    MULTS_3_13<=((others=> (others=>'0')));
    MULTS_3_14<=((others=> (others=>'0')));
    MULTS_3_15<=((others=> (others=>'0')));
    MULTS_3_16<=((others=> (others=>'0')));
    MULTS_3_17<=((others=> (others=>'0')));
    MULTS_3_18<=((others=> (others=>'0')));
    MULTS_3_19<=((others=> (others=>'0')));
    MULTS_3_20<=((others=> (others=>'0')));
    MULTS_3_21<=((others=> (others=>'0')));
    MULTS_3_22<=((others=> (others=>'0')));
    MULTS_3_23<=((others=> (others=>'0')));
    MULTS_3_24<=((others=> (others=>'0')));
    MULTS_3_25<=((others=> (others=>'0')));
    MULTS_3_26<=((others=> (others=>'0')));
    MULTS_3_27<=((others=> (others=>'0')));
    MULTS_3_28<=((others=> (others=>'0')));
    MULTS_3_29<=((others=> (others=>'0')));
    MULTS_3_30<=((others=> (others=>'0')));
    MULTS_3_31<=((others=> (others=>'0')));
    MULTS_3_32<=((others=> (others=>'0')));
    MULTS_3_33<=((others=> (others=>'0')));
    MULTS_3_34<=((others=> (others=>'0')));
    MULTS_3_35<=((others=> (others=>'0')));
    MULTS_3_36<=((others=> (others=>'0')));
    MULTS_3_37<=((others=> (others=>'0')));
    MULTS_3_38<=((others=> (others=>'0')));
    MULTS_3_39<=((others=> (others=>'0')));
    MULTS_3_40<=((others=> (others=>'0')));
    MULTS_3_41<=((others=> (others=>'0')));
    MULTS_3_42<=((others=> (others=>'0')));
    MULTS_3_43<=((others=> (others=>'0')));
    MULTS_3_44<=((others=> (others=>'0')));
    MULTS_3_45<=((others=> (others=>'0')));
    MULTS_3_46<=((others=> (others=>'0')));
    MULTS_3_47<=((others=> (others=>'0')));
    MULTS_3_48<=((others=> (others=>'0')));
    MULTS_3_49<=((others=> (others=>'0')));
    MULTS_3_50<=((others=> (others=>'0')));
    MULTS_3_51<=((others=> (others=>'0')));
    MULTS_3_52<=((others=> (others=>'0')));
    MULTS_3_53<=((others=> (others=>'0')));
    MULTS_3_54<=((others=> (others=>'0')));
    MULTS_3_55<=((others=> (others=>'0')));
    MULTS_3_56<=((others=> (others=>'0')));
    MULTS_3_57<=((others=> (others=>'0')));
    MULTS_3_58<=((others=> (others=>'0')));
    MULTS_3_59<=((others=> (others=>'0')));
    MULTS_3_60<=((others=> (others=>'0')));
    MULTS_3_61<=((others=> (others=>'0')));
    MULTS_3_62<=((others=> (others=>'0')));
    MULTS_3_63<=((others=> (others=>'0')));
    MULTS_3_64<=((others=> (others=>'0')));
    MULTS_3_65<=((others=> (others=>'0')));
    MULTS_3_66<=((others=> (others=>'0')));
    MULTS_3_67<=((others=> (others=>'0')));
    MULTS_3_68<=((others=> (others=>'0')));
    MULTS_3_69<=((others=> (others=>'0')));
    MULTS_3_70<=((others=> (others=>'0')));
    MULTS_3_71<=((others=> (others=>'0')));
    MULTS_3_72<=((others=> (others=>'0')));
    MULTS_3_73<=((others=> (others=>'0')));
    MULTS_3_74<=((others=> (others=>'0')));
    MULTS_3_75<=((others=> (others=>'0')));
    MULTS_3_76<=((others=> (others=>'0')));
    MULTS_3_77<=((others=> (others=>'0')));
    MULTS_3_78<=((others=> (others=>'0')));
    MULTS_3_79<=((others=> (others=>'0')));
    MULTS_3_80<=((others=> (others=>'0')));
    MULTS_3_81<=((others=> (others=>'0')));
    MULTS_3_82<=((others=> (others=>'0')));
    MULTS_3_83<=((others=> (others=>'0')));
    MULTS_3_84<=((others=> (others=>'0')));
    EN_SUM_MULT_4<='0';
    MULTS_4_1<=((others=> (others=>'0')));
    MULTS_4_2<=((others=> (others=>'0')));
    MULTS_4_3<=((others=> (others=>'0')));
    MULTS_4_4<=((others=> (others=>'0')));
    MULTS_4_5<=((others=> (others=>'0')));
    MULTS_4_6<=((others=> (others=>'0')));
    MULTS_4_7<=((others=> (others=>'0')));
    MULTS_4_8<=((others=> (others=>'0')));
    MULTS_4_9<=((others=> (others=>'0')));
    MULTS_4_10<=((others=> (others=>'0')));
    MULTS_4_11<=((others=> (others=>'0')));
    MULTS_4_12<=((others=> (others=>'0')));
    MULTS_4_13<=((others=> (others=>'0')));
    MULTS_4_14<=((others=> (others=>'0')));
    MULTS_4_15<=((others=> (others=>'0')));
    MULTS_4_16<=((others=> (others=>'0')));
    MULTS_4_17<=((others=> (others=>'0')));
    MULTS_4_18<=((others=> (others=>'0')));
    MULTS_4_19<=((others=> (others=>'0')));
    MULTS_4_20<=((others=> (others=>'0')));
    MULTS_4_21<=((others=> (others=>'0')));
    MULTS_4_22<=((others=> (others=>'0')));
    MULTS_4_23<=((others=> (others=>'0')));
    MULTS_4_24<=((others=> (others=>'0')));
    MULTS_4_25<=((others=> (others=>'0')));
    MULTS_4_26<=((others=> (others=>'0')));
    MULTS_4_27<=((others=> (others=>'0')));
    MULTS_4_28<=((others=> (others=>'0')));
    MULTS_4_29<=((others=> (others=>'0')));
    MULTS_4_30<=((others=> (others=>'0')));
    MULTS_4_31<=((others=> (others=>'0')));
    MULTS_4_32<=((others=> (others=>'0')));
    MULTS_4_33<=((others=> (others=>'0')));
    MULTS_4_34<=((others=> (others=>'0')));
    MULTS_4_35<=((others=> (others=>'0')));
    MULTS_4_36<=((others=> (others=>'0')));
    MULTS_4_37<=((others=> (others=>'0')));
    MULTS_4_38<=((others=> (others=>'0')));
    MULTS_4_39<=((others=> (others=>'0')));
    MULTS_4_40<=((others=> (others=>'0')));
    MULTS_4_41<=((others=> (others=>'0')));
    MULTS_4_42<=((others=> (others=>'0')));
    MULTS_4_43<=((others=> (others=>'0')));
    MULTS_4_44<=((others=> (others=>'0')));
    MULTS_4_45<=((others=> (others=>'0')));
    MULTS_4_46<=((others=> (others=>'0')));
    MULTS_4_47<=((others=> (others=>'0')));
    MULTS_4_48<=((others=> (others=>'0')));
    MULTS_4_49<=((others=> (others=>'0')));
    MULTS_4_50<=((others=> (others=>'0')));
    MULTS_4_51<=((others=> (others=>'0')));
    MULTS_4_52<=((others=> (others=>'0')));
    MULTS_4_53<=((others=> (others=>'0')));
    MULTS_4_54<=((others=> (others=>'0')));
    MULTS_4_55<=((others=> (others=>'0')));
    MULTS_4_56<=((others=> (others=>'0')));
    MULTS_4_57<=((others=> (others=>'0')));
    MULTS_4_58<=((others=> (others=>'0')));
    MULTS_4_59<=((others=> (others=>'0')));
    MULTS_4_60<=((others=> (others=>'0')));
    MULTS_4_61<=((others=> (others=>'0')));
    MULTS_4_62<=((others=> (others=>'0')));
    MULTS_4_63<=((others=> (others=>'0')));
    MULTS_4_64<=((others=> (others=>'0')));
    MULTS_4_65<=((others=> (others=>'0')));
    MULTS_4_66<=((others=> (others=>'0')));
    MULTS_4_67<=((others=> (others=>'0')));
    MULTS_4_68<=((others=> (others=>'0')));
    MULTS_4_69<=((others=> (others=>'0')));
    MULTS_4_70<=((others=> (others=>'0')));
    MULTS_4_71<=((others=> (others=>'0')));
    MULTS_4_72<=((others=> (others=>'0')));
    MULTS_4_73<=((others=> (others=>'0')));
    MULTS_4_74<=((others=> (others=>'0')));
    MULTS_4_75<=((others=> (others=>'0')));
    MULTS_4_76<=((others=> (others=>'0')));
    MULTS_4_77<=((others=> (others=>'0')));
    MULTS_4_78<=((others=> (others=>'0')));
    MULTS_4_79<=((others=> (others=>'0')));
    MULTS_4_80<=((others=> (others=>'0')));
    MULTS_4_81<=((others=> (others=>'0')));
    MULTS_4_82<=((others=> (others=>'0')));
    MULTS_4_83<=((others=> (others=>'0')));
    MULTS_4_84<=((others=> (others=>'0')));
    EN_SUM_MULT_5<='0';
    MULTS_5_1<=((others=> (others=>'0')));
    MULTS_5_2<=((others=> (others=>'0')));
    MULTS_5_3<=((others=> (others=>'0')));
    MULTS_5_4<=((others=> (others=>'0')));
    MULTS_5_5<=((others=> (others=>'0')));
    MULTS_5_6<=((others=> (others=>'0')));
    MULTS_5_7<=((others=> (others=>'0')));
    MULTS_5_8<=((others=> (others=>'0')));
    MULTS_5_9<=((others=> (others=>'0')));
    MULTS_5_10<=((others=> (others=>'0')));
    MULTS_5_11<=((others=> (others=>'0')));
    MULTS_5_12<=((others=> (others=>'0')));
    MULTS_5_13<=((others=> (others=>'0')));
    MULTS_5_14<=((others=> (others=>'0')));
    MULTS_5_15<=((others=> (others=>'0')));
    MULTS_5_16<=((others=> (others=>'0')));
    MULTS_5_17<=((others=> (others=>'0')));
    MULTS_5_18<=((others=> (others=>'0')));
    MULTS_5_19<=((others=> (others=>'0')));
    MULTS_5_20<=((others=> (others=>'0')));
    MULTS_5_21<=((others=> (others=>'0')));
    MULTS_5_22<=((others=> (others=>'0')));
    MULTS_5_23<=((others=> (others=>'0')));
    MULTS_5_24<=((others=> (others=>'0')));
    MULTS_5_25<=((others=> (others=>'0')));
    MULTS_5_26<=((others=> (others=>'0')));
    MULTS_5_27<=((others=> (others=>'0')));
    MULTS_5_28<=((others=> (others=>'0')));
    MULTS_5_29<=((others=> (others=>'0')));
    MULTS_5_30<=((others=> (others=>'0')));
    MULTS_5_31<=((others=> (others=>'0')));
    MULTS_5_32<=((others=> (others=>'0')));
    MULTS_5_33<=((others=> (others=>'0')));
    MULTS_5_34<=((others=> (others=>'0')));
    MULTS_5_35<=((others=> (others=>'0')));
    MULTS_5_36<=((others=> (others=>'0')));
    MULTS_5_37<=((others=> (others=>'0')));
    MULTS_5_38<=((others=> (others=>'0')));
    MULTS_5_39<=((others=> (others=>'0')));
    MULTS_5_40<=((others=> (others=>'0')));
    MULTS_5_41<=((others=> (others=>'0')));
    MULTS_5_42<=((others=> (others=>'0')));
    MULTS_5_43<=((others=> (others=>'0')));
    MULTS_5_44<=((others=> (others=>'0')));
    MULTS_5_45<=((others=> (others=>'0')));
    MULTS_5_46<=((others=> (others=>'0')));
    MULTS_5_47<=((others=> (others=>'0')));
    MULTS_5_48<=((others=> (others=>'0')));
    MULTS_5_49<=((others=> (others=>'0')));
    MULTS_5_50<=((others=> (others=>'0')));
    MULTS_5_51<=((others=> (others=>'0')));
    MULTS_5_52<=((others=> (others=>'0')));
    MULTS_5_53<=((others=> (others=>'0')));
    MULTS_5_54<=((others=> (others=>'0')));
    MULTS_5_55<=((others=> (others=>'0')));
    MULTS_5_56<=((others=> (others=>'0')));
    MULTS_5_57<=((others=> (others=>'0')));
    MULTS_5_58<=((others=> (others=>'0')));
    MULTS_5_59<=((others=> (others=>'0')));
    MULTS_5_60<=((others=> (others=>'0')));
    MULTS_5_61<=((others=> (others=>'0')));
    MULTS_5_62<=((others=> (others=>'0')));
    MULTS_5_63<=((others=> (others=>'0')));
    MULTS_5_64<=((others=> (others=>'0')));
    MULTS_5_65<=((others=> (others=>'0')));
    MULTS_5_66<=((others=> (others=>'0')));
    MULTS_5_67<=((others=> (others=>'0')));
    MULTS_5_68<=((others=> (others=>'0')));
    MULTS_5_69<=((others=> (others=>'0')));
    MULTS_5_70<=((others=> (others=>'0')));
    MULTS_5_71<=((others=> (others=>'0')));
    MULTS_5_72<=((others=> (others=>'0')));
    MULTS_5_73<=((others=> (others=>'0')));
    MULTS_5_74<=((others=> (others=>'0')));
    MULTS_5_75<=((others=> (others=>'0')));
    MULTS_5_76<=((others=> (others=>'0')));
    MULTS_5_77<=((others=> (others=>'0')));
    MULTS_5_78<=((others=> (others=>'0')));
    MULTS_5_79<=((others=> (others=>'0')));
    MULTS_5_80<=((others=> (others=>'0')));
    MULTS_5_81<=((others=> (others=>'0')));
    MULTS_5_82<=((others=> (others=>'0')));
    MULTS_5_83<=((others=> (others=>'0')));
    MULTS_5_84<=((others=> (others=>'0')));
    EN_SUM_MULT_6<='0';
    MULTS_6_1<=((others=> (others=>'0')));
    MULTS_6_2<=((others=> (others=>'0')));
    MULTS_6_3<=((others=> (others=>'0')));
    MULTS_6_4<=((others=> (others=>'0')));
    MULTS_6_5<=((others=> (others=>'0')));
    MULTS_6_6<=((others=> (others=>'0')));
    MULTS_6_7<=((others=> (others=>'0')));
    MULTS_6_8<=((others=> (others=>'0')));
    MULTS_6_9<=((others=> (others=>'0')));
    MULTS_6_10<=((others=> (others=>'0')));
    MULTS_6_11<=((others=> (others=>'0')));
    MULTS_6_12<=((others=> (others=>'0')));
    MULTS_6_13<=((others=> (others=>'0')));
    MULTS_6_14<=((others=> (others=>'0')));
    MULTS_6_15<=((others=> (others=>'0')));
    MULTS_6_16<=((others=> (others=>'0')));
    MULTS_6_17<=((others=> (others=>'0')));
    MULTS_6_18<=((others=> (others=>'0')));
    MULTS_6_19<=((others=> (others=>'0')));
    MULTS_6_20<=((others=> (others=>'0')));
    MULTS_6_21<=((others=> (others=>'0')));
    MULTS_6_22<=((others=> (others=>'0')));
    MULTS_6_23<=((others=> (others=>'0')));
    MULTS_6_24<=((others=> (others=>'0')));
    MULTS_6_25<=((others=> (others=>'0')));
    MULTS_6_26<=((others=> (others=>'0')));
    MULTS_6_27<=((others=> (others=>'0')));
    MULTS_6_28<=((others=> (others=>'0')));
    MULTS_6_29<=((others=> (others=>'0')));
    MULTS_6_30<=((others=> (others=>'0')));
    MULTS_6_31<=((others=> (others=>'0')));
    MULTS_6_32<=((others=> (others=>'0')));
    MULTS_6_33<=((others=> (others=>'0')));
    MULTS_6_34<=((others=> (others=>'0')));
    MULTS_6_35<=((others=> (others=>'0')));
    MULTS_6_36<=((others=> (others=>'0')));
    MULTS_6_37<=((others=> (others=>'0')));
    MULTS_6_38<=((others=> (others=>'0')));
    MULTS_6_39<=((others=> (others=>'0')));
    MULTS_6_40<=((others=> (others=>'0')));
    MULTS_6_41<=((others=> (others=>'0')));
    MULTS_6_42<=((others=> (others=>'0')));
    MULTS_6_43<=((others=> (others=>'0')));
    MULTS_6_44<=((others=> (others=>'0')));
    MULTS_6_45<=((others=> (others=>'0')));
    MULTS_6_46<=((others=> (others=>'0')));
    MULTS_6_47<=((others=> (others=>'0')));
    MULTS_6_48<=((others=> (others=>'0')));
    MULTS_6_49<=((others=> (others=>'0')));
    MULTS_6_50<=((others=> (others=>'0')));
    MULTS_6_51<=((others=> (others=>'0')));
    MULTS_6_52<=((others=> (others=>'0')));
    MULTS_6_53<=((others=> (others=>'0')));
    MULTS_6_54<=((others=> (others=>'0')));
    MULTS_6_55<=((others=> (others=>'0')));
    MULTS_6_56<=((others=> (others=>'0')));
    MULTS_6_57<=((others=> (others=>'0')));
    MULTS_6_58<=((others=> (others=>'0')));
    MULTS_6_59<=((others=> (others=>'0')));
    MULTS_6_60<=((others=> (others=>'0')));
    MULTS_6_61<=((others=> (others=>'0')));
    MULTS_6_62<=((others=> (others=>'0')));
    MULTS_6_63<=((others=> (others=>'0')));
    MULTS_6_64<=((others=> (others=>'0')));
    MULTS_6_65<=((others=> (others=>'0')));
    MULTS_6_66<=((others=> (others=>'0')));
    MULTS_6_67<=((others=> (others=>'0')));
    MULTS_6_68<=((others=> (others=>'0')));
    MULTS_6_69<=((others=> (others=>'0')));
    MULTS_6_70<=((others=> (others=>'0')));
    MULTS_6_71<=((others=> (others=>'0')));
    MULTS_6_72<=((others=> (others=>'0')));
    MULTS_6_73<=((others=> (others=>'0')));
    MULTS_6_74<=((others=> (others=>'0')));
    MULTS_6_75<=((others=> (others=>'0')));
    MULTS_6_76<=((others=> (others=>'0')));
    MULTS_6_77<=((others=> (others=>'0')));
    MULTS_6_78<=((others=> (others=>'0')));
    MULTS_6_79<=((others=> (others=>'0')));
    MULTS_6_80<=((others=> (others=>'0')));
    MULTS_6_81<=((others=> (others=>'0')));
    MULTS_6_82<=((others=> (others=>'0')));
    MULTS_6_83<=((others=> (others=>'0')));
    MULTS_6_84<=((others=> (others=>'0')));
    EN_SUM_MULT_7<='0';
    MULTS_7_1<=((others=> (others=>'0')));
    MULTS_7_2<=((others=> (others=>'0')));
    MULTS_7_3<=((others=> (others=>'0')));
    MULTS_7_4<=((others=> (others=>'0')));
    MULTS_7_5<=((others=> (others=>'0')));
    MULTS_7_6<=((others=> (others=>'0')));
    MULTS_7_7<=((others=> (others=>'0')));
    MULTS_7_8<=((others=> (others=>'0')));
    MULTS_7_9<=((others=> (others=>'0')));
    MULTS_7_10<=((others=> (others=>'0')));
    MULTS_7_11<=((others=> (others=>'0')));
    MULTS_7_12<=((others=> (others=>'0')));
    MULTS_7_13<=((others=> (others=>'0')));
    MULTS_7_14<=((others=> (others=>'0')));
    MULTS_7_15<=((others=> (others=>'0')));
    MULTS_7_16<=((others=> (others=>'0')));
    MULTS_7_17<=((others=> (others=>'0')));
    MULTS_7_18<=((others=> (others=>'0')));
    MULTS_7_19<=((others=> (others=>'0')));
    MULTS_7_20<=((others=> (others=>'0')));
    MULTS_7_21<=((others=> (others=>'0')));
    MULTS_7_22<=((others=> (others=>'0')));
    MULTS_7_23<=((others=> (others=>'0')));
    MULTS_7_24<=((others=> (others=>'0')));
    MULTS_7_25<=((others=> (others=>'0')));
    MULTS_7_26<=((others=> (others=>'0')));
    MULTS_7_27<=((others=> (others=>'0')));
    MULTS_7_28<=((others=> (others=>'0')));
    MULTS_7_29<=((others=> (others=>'0')));
    MULTS_7_30<=((others=> (others=>'0')));
    MULTS_7_31<=((others=> (others=>'0')));
    MULTS_7_32<=((others=> (others=>'0')));
    MULTS_7_33<=((others=> (others=>'0')));
    MULTS_7_34<=((others=> (others=>'0')));
    MULTS_7_35<=((others=> (others=>'0')));
    MULTS_7_36<=((others=> (others=>'0')));
    MULTS_7_37<=((others=> (others=>'0')));
    MULTS_7_38<=((others=> (others=>'0')));
    MULTS_7_39<=((others=> (others=>'0')));
    MULTS_7_40<=((others=> (others=>'0')));
    MULTS_7_41<=((others=> (others=>'0')));
    MULTS_7_42<=((others=> (others=>'0')));
    MULTS_7_43<=((others=> (others=>'0')));
    MULTS_7_44<=((others=> (others=>'0')));
    MULTS_7_45<=((others=> (others=>'0')));
    MULTS_7_46<=((others=> (others=>'0')));
    MULTS_7_47<=((others=> (others=>'0')));
    MULTS_7_48<=((others=> (others=>'0')));
    MULTS_7_49<=((others=> (others=>'0')));
    MULTS_7_50<=((others=> (others=>'0')));
    MULTS_7_51<=((others=> (others=>'0')));
    MULTS_7_52<=((others=> (others=>'0')));
    MULTS_7_53<=((others=> (others=>'0')));
    MULTS_7_54<=((others=> (others=>'0')));
    MULTS_7_55<=((others=> (others=>'0')));
    MULTS_7_56<=((others=> (others=>'0')));
    MULTS_7_57<=((others=> (others=>'0')));
    MULTS_7_58<=((others=> (others=>'0')));
    MULTS_7_59<=((others=> (others=>'0')));
    MULTS_7_60<=((others=> (others=>'0')));
    MULTS_7_61<=((others=> (others=>'0')));
    MULTS_7_62<=((others=> (others=>'0')));
    MULTS_7_63<=((others=> (others=>'0')));
    MULTS_7_64<=((others=> (others=>'0')));
    MULTS_7_65<=((others=> (others=>'0')));
    MULTS_7_66<=((others=> (others=>'0')));
    MULTS_7_67<=((others=> (others=>'0')));
    MULTS_7_68<=((others=> (others=>'0')));
    MULTS_7_69<=((others=> (others=>'0')));
    MULTS_7_70<=((others=> (others=>'0')));
    MULTS_7_71<=((others=> (others=>'0')));
    MULTS_7_72<=((others=> (others=>'0')));
    MULTS_7_73<=((others=> (others=>'0')));
    MULTS_7_74<=((others=> (others=>'0')));
    MULTS_7_75<=((others=> (others=>'0')));
    MULTS_7_76<=((others=> (others=>'0')));
    MULTS_7_77<=((others=> (others=>'0')));
    MULTS_7_78<=((others=> (others=>'0')));
    MULTS_7_79<=((others=> (others=>'0')));
    MULTS_7_80<=((others=> (others=>'0')));
    MULTS_7_81<=((others=> (others=>'0')));
    MULTS_7_82<=((others=> (others=>'0')));
    MULTS_7_83<=((others=> (others=>'0')));
    MULTS_7_84<=((others=> (others=>'0')));

------------------------------------------------ PROCESS START------------------------------------------------------
	  
   else 	
	if EN_LOC_STREAM_8='1' and EN_STREAM= '1' and OUT_PIXEL_COUNT<VALID_CYCLES  then    -- check valid data and enable stream
		
		if  FRST_TIM_EN_8='1' then EN_NXT_LYR_8<='1';end if;

			MULT_1(0)<=signed(DIN_1_8)*signed(FMAP_1_1);
			MULT_2(0)<=signed(DIN_2_8)*signed(FMAP_1_2);
			MULT_3(0)<=signed(DIN_3_8)*signed(FMAP_1_3);
			MULT_4(0)<=signed(DIN_4_8)*signed(FMAP_1_4);
			MULT_5(0)<=signed(DIN_5_8)*signed(FMAP_1_5);
			MULT_6(0)<=signed(DIN_6_8)*signed(FMAP_1_6);
			MULT_7(0)<=signed(DIN_7_8)*signed(FMAP_1_7);
			MULT_8(0)<=signed(DIN_8_8)*signed(FMAP_1_8);
			MULT_9(0)<=signed(DIN_9_8)*signed(FMAP_1_9);
			MULT_10(0)<=signed(DIN_10_8)*signed(FMAP_1_10);
			MULT_11(0)<=signed(DIN_11_8)*signed(FMAP_1_11);
			MULT_12(0)<=signed(DIN_12_8)*signed(FMAP_1_12);
			MULT_13(0)<=signed(DIN_13_8)*signed(FMAP_1_13);
			MULT_14(0)<=signed(DIN_14_8)*signed(FMAP_1_14);
			MULT_15(0)<=signed(DIN_15_8)*signed(FMAP_1_15);
			MULT_16(0)<=signed(DIN_16_8)*signed(FMAP_1_16);
			MULT_17(0)<=signed(DIN_17_8)*signed(FMAP_1_17);
			MULT_18(0)<=signed(DIN_18_8)*signed(FMAP_1_18);
			MULT_19(0)<=signed(DIN_19_8)*signed(FMAP_1_19);
			MULT_20(0)<=signed(DIN_20_8)*signed(FMAP_1_20);
			MULT_21(0)<=signed(DIN_21_8)*signed(FMAP_1_21);
			MULT_22(0)<=signed(DIN_22_8)*signed(FMAP_1_22);
			MULT_23(0)<=signed(DIN_23_8)*signed(FMAP_1_23);
			MULT_24(0)<=signed(DIN_24_8)*signed(FMAP_1_24);
			MULT_25(0)<=signed(DIN_25_8)*signed(FMAP_1_25);
			MULT_26(0)<=signed(DIN_26_8)*signed(FMAP_1_26);
			MULT_27(0)<=signed(DIN_27_8)*signed(FMAP_1_27);
			MULT_28(0)<=signed(DIN_28_8)*signed(FMAP_1_28);
			MULT_29(0)<=signed(DIN_29_8)*signed(FMAP_1_29);
			MULT_30(0)<=signed(DIN_30_8)*signed(FMAP_1_30);
			MULT_31(0)<=signed(DIN_31_8)*signed(FMAP_1_31);
			MULT_32(0)<=signed(DIN_32_8)*signed(FMAP_1_32);
			MULT_33(0)<=signed(DIN_33_8)*signed(FMAP_1_33);
			MULT_34(0)<=signed(DIN_34_8)*signed(FMAP_1_34);
			MULT_35(0)<=signed(DIN_35_8)*signed(FMAP_1_35);
			MULT_36(0)<=signed(DIN_36_8)*signed(FMAP_1_36);
			MULT_37(0)<=signed(DIN_37_8)*signed(FMAP_1_37);
			MULT_38(0)<=signed(DIN_38_8)*signed(FMAP_1_38);
			MULT_39(0)<=signed(DIN_39_8)*signed(FMAP_1_39);
			MULT_40(0)<=signed(DIN_40_8)*signed(FMAP_1_40);
			MULT_41(0)<=signed(DIN_41_8)*signed(FMAP_1_41);
			MULT_42(0)<=signed(DIN_42_8)*signed(FMAP_1_42);
			MULT_43(0)<=signed(DIN_43_8)*signed(FMAP_1_43);
			MULT_44(0)<=signed(DIN_44_8)*signed(FMAP_1_44);
			MULT_45(0)<=signed(DIN_45_8)*signed(FMAP_1_45);
			MULT_46(0)<=signed(DIN_46_8)*signed(FMAP_1_46);
			MULT_47(0)<=signed(DIN_47_8)*signed(FMAP_1_47);
			MULT_48(0)<=signed(DIN_48_8)*signed(FMAP_1_48);
			MULT_49(0)<=signed(DIN_49_8)*signed(FMAP_1_49);
			MULT_50(0)<=signed(DIN_50_8)*signed(FMAP_1_50);
			MULT_51(0)<=signed(DIN_51_8)*signed(FMAP_1_51);
			MULT_52(0)<=signed(DIN_52_8)*signed(FMAP_1_52);
			MULT_53(0)<=signed(DIN_53_8)*signed(FMAP_1_53);
			MULT_54(0)<=signed(DIN_54_8)*signed(FMAP_1_54);
			MULT_55(0)<=signed(DIN_55_8)*signed(FMAP_1_55);
			MULT_56(0)<=signed(DIN_56_8)*signed(FMAP_1_56);
			MULT_57(0)<=signed(DIN_57_8)*signed(FMAP_1_57);
			MULT_58(0)<=signed(DIN_58_8)*signed(FMAP_1_58);
			MULT_59(0)<=signed(DIN_59_8)*signed(FMAP_1_59);
			MULT_60(0)<=signed(DIN_60_8)*signed(FMAP_1_60);
			MULT_61(0)<=signed(DIN_61_8)*signed(FMAP_1_61);
			MULT_62(0)<=signed(DIN_62_8)*signed(FMAP_1_62);
			MULT_63(0)<=signed(DIN_63_8)*signed(FMAP_1_63);
			MULT_64(0)<=signed(DIN_64_8)*signed(FMAP_1_64);
			MULT_65(0)<=signed(DIN_65_8)*signed(FMAP_1_65);
			MULT_66(0)<=signed(DIN_66_8)*signed(FMAP_1_66);
			MULT_67(0)<=signed(DIN_67_8)*signed(FMAP_1_67);
			MULT_68(0)<=signed(DIN_68_8)*signed(FMAP_1_68);
			MULT_69(0)<=signed(DIN_69_8)*signed(FMAP_1_69);
			MULT_70(0)<=signed(DIN_70_8)*signed(FMAP_1_70);
			MULT_71(0)<=signed(DIN_71_8)*signed(FMAP_1_71);
			MULT_72(0)<=signed(DIN_72_8)*signed(FMAP_1_72);
			MULT_73(0)<=signed(DIN_73_8)*signed(FMAP_1_73);
			MULT_74(0)<=signed(DIN_74_8)*signed(FMAP_1_74);
			MULT_75(0)<=signed(DIN_75_8)*signed(FMAP_1_75);
			MULT_76(0)<=signed(DIN_76_8)*signed(FMAP_1_76);
			MULT_77(0)<=signed(DIN_77_8)*signed(FMAP_1_77);
			MULT_78(0)<=signed(DIN_78_8)*signed(FMAP_1_78);
			MULT_79(0)<=signed(DIN_79_8)*signed(FMAP_1_79);
			MULT_80(0)<=signed(DIN_80_8)*signed(FMAP_1_80);
			MULT_81(0)<=signed(DIN_81_8)*signed(FMAP_1_81);
			MULT_82(0)<=signed(DIN_82_8)*signed(FMAP_1_82);
			MULT_83(0)<=signed(DIN_83_8)*signed(FMAP_1_83);
			MULT_84(0)<=signed(DIN_84_8)*signed(FMAP_1_84);

			MULT_1(1)<=signed(DIN_1_8)*signed(FMAP_2_1);
			MULT_2(1)<=signed(DIN_2_8)*signed(FMAP_2_2);
			MULT_3(1)<=signed(DIN_3_8)*signed(FMAP_2_3);
			MULT_4(1)<=signed(DIN_4_8)*signed(FMAP_2_4);
			MULT_5(1)<=signed(DIN_5_8)*signed(FMAP_2_5);
			MULT_6(1)<=signed(DIN_6_8)*signed(FMAP_2_6);
			MULT_7(1)<=signed(DIN_7_8)*signed(FMAP_2_7);
			MULT_8(1)<=signed(DIN_8_8)*signed(FMAP_2_8);
			MULT_9(1)<=signed(DIN_9_8)*signed(FMAP_2_9);
			MULT_10(1)<=signed(DIN_10_8)*signed(FMAP_2_10);
			MULT_11(1)<=signed(DIN_11_8)*signed(FMAP_2_11);
			MULT_12(1)<=signed(DIN_12_8)*signed(FMAP_2_12);
			MULT_13(1)<=signed(DIN_13_8)*signed(FMAP_2_13);
			MULT_14(1)<=signed(DIN_14_8)*signed(FMAP_2_14);
			MULT_15(1)<=signed(DIN_15_8)*signed(FMAP_2_15);
			MULT_16(1)<=signed(DIN_16_8)*signed(FMAP_2_16);
			MULT_17(1)<=signed(DIN_17_8)*signed(FMAP_2_17);
			MULT_18(1)<=signed(DIN_18_8)*signed(FMAP_2_18);
			MULT_19(1)<=signed(DIN_19_8)*signed(FMAP_2_19);
			MULT_20(1)<=signed(DIN_20_8)*signed(FMAP_2_20);
			MULT_21(1)<=signed(DIN_21_8)*signed(FMAP_2_21);
			MULT_22(1)<=signed(DIN_22_8)*signed(FMAP_2_22);
			MULT_23(1)<=signed(DIN_23_8)*signed(FMAP_2_23);
			MULT_24(1)<=signed(DIN_24_8)*signed(FMAP_2_24);
			MULT_25(1)<=signed(DIN_25_8)*signed(FMAP_2_25);
			MULT_26(1)<=signed(DIN_26_8)*signed(FMAP_2_26);
			MULT_27(1)<=signed(DIN_27_8)*signed(FMAP_2_27);
			MULT_28(1)<=signed(DIN_28_8)*signed(FMAP_2_28);
			MULT_29(1)<=signed(DIN_29_8)*signed(FMAP_2_29);
			MULT_30(1)<=signed(DIN_30_8)*signed(FMAP_2_30);
			MULT_31(1)<=signed(DIN_31_8)*signed(FMAP_2_31);
			MULT_32(1)<=signed(DIN_32_8)*signed(FMAP_2_32);
			MULT_33(1)<=signed(DIN_33_8)*signed(FMAP_2_33);
			MULT_34(1)<=signed(DIN_34_8)*signed(FMAP_2_34);
			MULT_35(1)<=signed(DIN_35_8)*signed(FMAP_2_35);
			MULT_36(1)<=signed(DIN_36_8)*signed(FMAP_2_36);
			MULT_37(1)<=signed(DIN_37_8)*signed(FMAP_2_37);
			MULT_38(1)<=signed(DIN_38_8)*signed(FMAP_2_38);
			MULT_39(1)<=signed(DIN_39_8)*signed(FMAP_2_39);
			MULT_40(1)<=signed(DIN_40_8)*signed(FMAP_2_40);
			MULT_41(1)<=signed(DIN_41_8)*signed(FMAP_2_41);
			MULT_42(1)<=signed(DIN_42_8)*signed(FMAP_2_42);
			MULT_43(1)<=signed(DIN_43_8)*signed(FMAP_2_43);
			MULT_44(1)<=signed(DIN_44_8)*signed(FMAP_2_44);
			MULT_45(1)<=signed(DIN_45_8)*signed(FMAP_2_45);
			MULT_46(1)<=signed(DIN_46_8)*signed(FMAP_2_46);
			MULT_47(1)<=signed(DIN_47_8)*signed(FMAP_2_47);
			MULT_48(1)<=signed(DIN_48_8)*signed(FMAP_2_48);
			MULT_49(1)<=signed(DIN_49_8)*signed(FMAP_2_49);
			MULT_50(1)<=signed(DIN_50_8)*signed(FMAP_2_50);
			MULT_51(1)<=signed(DIN_51_8)*signed(FMAP_2_51);
			MULT_52(1)<=signed(DIN_52_8)*signed(FMAP_2_52);
			MULT_53(1)<=signed(DIN_53_8)*signed(FMAP_2_53);
			MULT_54(1)<=signed(DIN_54_8)*signed(FMAP_2_54);
			MULT_55(1)<=signed(DIN_55_8)*signed(FMAP_2_55);
			MULT_56(1)<=signed(DIN_56_8)*signed(FMAP_2_56);
			MULT_57(1)<=signed(DIN_57_8)*signed(FMAP_2_57);
			MULT_58(1)<=signed(DIN_58_8)*signed(FMAP_2_58);
			MULT_59(1)<=signed(DIN_59_8)*signed(FMAP_2_59);
			MULT_60(1)<=signed(DIN_60_8)*signed(FMAP_2_60);
			MULT_61(1)<=signed(DIN_61_8)*signed(FMAP_2_61);
			MULT_62(1)<=signed(DIN_62_8)*signed(FMAP_2_62);
			MULT_63(1)<=signed(DIN_63_8)*signed(FMAP_2_63);
			MULT_64(1)<=signed(DIN_64_8)*signed(FMAP_2_64);
			MULT_65(1)<=signed(DIN_65_8)*signed(FMAP_2_65);
			MULT_66(1)<=signed(DIN_66_8)*signed(FMAP_2_66);
			MULT_67(1)<=signed(DIN_67_8)*signed(FMAP_2_67);
			MULT_68(1)<=signed(DIN_68_8)*signed(FMAP_2_68);
			MULT_69(1)<=signed(DIN_69_8)*signed(FMAP_2_69);
			MULT_70(1)<=signed(DIN_70_8)*signed(FMAP_2_70);
			MULT_71(1)<=signed(DIN_71_8)*signed(FMAP_2_71);
			MULT_72(1)<=signed(DIN_72_8)*signed(FMAP_2_72);
			MULT_73(1)<=signed(DIN_73_8)*signed(FMAP_2_73);
			MULT_74(1)<=signed(DIN_74_8)*signed(FMAP_2_74);
			MULT_75(1)<=signed(DIN_75_8)*signed(FMAP_2_75);
			MULT_76(1)<=signed(DIN_76_8)*signed(FMAP_2_76);
			MULT_77(1)<=signed(DIN_77_8)*signed(FMAP_2_77);
			MULT_78(1)<=signed(DIN_78_8)*signed(FMAP_2_78);
			MULT_79(1)<=signed(DIN_79_8)*signed(FMAP_2_79);
			MULT_80(1)<=signed(DIN_80_8)*signed(FMAP_2_80);
			MULT_81(1)<=signed(DIN_81_8)*signed(FMAP_2_81);
			MULT_82(1)<=signed(DIN_82_8)*signed(FMAP_2_82);
			MULT_83(1)<=signed(DIN_83_8)*signed(FMAP_2_83);
			MULT_84(1)<=signed(DIN_84_8)*signed(FMAP_2_84);

			MULT_1(2)<=signed(DIN_1_8)*signed(FMAP_3_1);
			MULT_2(2)<=signed(DIN_2_8)*signed(FMAP_3_2);
			MULT_3(2)<=signed(DIN_3_8)*signed(FMAP_3_3);
			MULT_4(2)<=signed(DIN_4_8)*signed(FMAP_3_4);
			MULT_5(2)<=signed(DIN_5_8)*signed(FMAP_3_5);
			MULT_6(2)<=signed(DIN_6_8)*signed(FMAP_3_6);
			MULT_7(2)<=signed(DIN_7_8)*signed(FMAP_3_7);
			MULT_8(2)<=signed(DIN_8_8)*signed(FMAP_3_8);
			MULT_9(2)<=signed(DIN_9_8)*signed(FMAP_3_9);
			MULT_10(2)<=signed(DIN_10_8)*signed(FMAP_3_10);
			MULT_11(2)<=signed(DIN_11_8)*signed(FMAP_3_11);
			MULT_12(2)<=signed(DIN_12_8)*signed(FMAP_3_12);
			MULT_13(2)<=signed(DIN_13_8)*signed(FMAP_3_13);
			MULT_14(2)<=signed(DIN_14_8)*signed(FMAP_3_14);
			MULT_15(2)<=signed(DIN_15_8)*signed(FMAP_3_15);
			MULT_16(2)<=signed(DIN_16_8)*signed(FMAP_3_16);
			MULT_17(2)<=signed(DIN_17_8)*signed(FMAP_3_17);
			MULT_18(2)<=signed(DIN_18_8)*signed(FMAP_3_18);
			MULT_19(2)<=signed(DIN_19_8)*signed(FMAP_3_19);
			MULT_20(2)<=signed(DIN_20_8)*signed(FMAP_3_20);
			MULT_21(2)<=signed(DIN_21_8)*signed(FMAP_3_21);
			MULT_22(2)<=signed(DIN_22_8)*signed(FMAP_3_22);
			MULT_23(2)<=signed(DIN_23_8)*signed(FMAP_3_23);
			MULT_24(2)<=signed(DIN_24_8)*signed(FMAP_3_24);
			MULT_25(2)<=signed(DIN_25_8)*signed(FMAP_3_25);
			MULT_26(2)<=signed(DIN_26_8)*signed(FMAP_3_26);
			MULT_27(2)<=signed(DIN_27_8)*signed(FMAP_3_27);
			MULT_28(2)<=signed(DIN_28_8)*signed(FMAP_3_28);
			MULT_29(2)<=signed(DIN_29_8)*signed(FMAP_3_29);
			MULT_30(2)<=signed(DIN_30_8)*signed(FMAP_3_30);
			MULT_31(2)<=signed(DIN_31_8)*signed(FMAP_3_31);
			MULT_32(2)<=signed(DIN_32_8)*signed(FMAP_3_32);
			MULT_33(2)<=signed(DIN_33_8)*signed(FMAP_3_33);
			MULT_34(2)<=signed(DIN_34_8)*signed(FMAP_3_34);
			MULT_35(2)<=signed(DIN_35_8)*signed(FMAP_3_35);
			MULT_36(2)<=signed(DIN_36_8)*signed(FMAP_3_36);
			MULT_37(2)<=signed(DIN_37_8)*signed(FMAP_3_37);
			MULT_38(2)<=signed(DIN_38_8)*signed(FMAP_3_38);
			MULT_39(2)<=signed(DIN_39_8)*signed(FMAP_3_39);
			MULT_40(2)<=signed(DIN_40_8)*signed(FMAP_3_40);
			MULT_41(2)<=signed(DIN_41_8)*signed(FMAP_3_41);
			MULT_42(2)<=signed(DIN_42_8)*signed(FMAP_3_42);
			MULT_43(2)<=signed(DIN_43_8)*signed(FMAP_3_43);
			MULT_44(2)<=signed(DIN_44_8)*signed(FMAP_3_44);
			MULT_45(2)<=signed(DIN_45_8)*signed(FMAP_3_45);
			MULT_46(2)<=signed(DIN_46_8)*signed(FMAP_3_46);
			MULT_47(2)<=signed(DIN_47_8)*signed(FMAP_3_47);
			MULT_48(2)<=signed(DIN_48_8)*signed(FMAP_3_48);
			MULT_49(2)<=signed(DIN_49_8)*signed(FMAP_3_49);
			MULT_50(2)<=signed(DIN_50_8)*signed(FMAP_3_50);
			MULT_51(2)<=signed(DIN_51_8)*signed(FMAP_3_51);
			MULT_52(2)<=signed(DIN_52_8)*signed(FMAP_3_52);
			MULT_53(2)<=signed(DIN_53_8)*signed(FMAP_3_53);
			MULT_54(2)<=signed(DIN_54_8)*signed(FMAP_3_54);
			MULT_55(2)<=signed(DIN_55_8)*signed(FMAP_3_55);
			MULT_56(2)<=signed(DIN_56_8)*signed(FMAP_3_56);
			MULT_57(2)<=signed(DIN_57_8)*signed(FMAP_3_57);
			MULT_58(2)<=signed(DIN_58_8)*signed(FMAP_3_58);
			MULT_59(2)<=signed(DIN_59_8)*signed(FMAP_3_59);
			MULT_60(2)<=signed(DIN_60_8)*signed(FMAP_3_60);
			MULT_61(2)<=signed(DIN_61_8)*signed(FMAP_3_61);
			MULT_62(2)<=signed(DIN_62_8)*signed(FMAP_3_62);
			MULT_63(2)<=signed(DIN_63_8)*signed(FMAP_3_63);
			MULT_64(2)<=signed(DIN_64_8)*signed(FMAP_3_64);
			MULT_65(2)<=signed(DIN_65_8)*signed(FMAP_3_65);
			MULT_66(2)<=signed(DIN_66_8)*signed(FMAP_3_66);
			MULT_67(2)<=signed(DIN_67_8)*signed(FMAP_3_67);
			MULT_68(2)<=signed(DIN_68_8)*signed(FMAP_3_68);
			MULT_69(2)<=signed(DIN_69_8)*signed(FMAP_3_69);
			MULT_70(2)<=signed(DIN_70_8)*signed(FMAP_3_70);
			MULT_71(2)<=signed(DIN_71_8)*signed(FMAP_3_71);
			MULT_72(2)<=signed(DIN_72_8)*signed(FMAP_3_72);
			MULT_73(2)<=signed(DIN_73_8)*signed(FMAP_3_73);
			MULT_74(2)<=signed(DIN_74_8)*signed(FMAP_3_74);
			MULT_75(2)<=signed(DIN_75_8)*signed(FMAP_3_75);
			MULT_76(2)<=signed(DIN_76_8)*signed(FMAP_3_76);
			MULT_77(2)<=signed(DIN_77_8)*signed(FMAP_3_77);
			MULT_78(2)<=signed(DIN_78_8)*signed(FMAP_3_78);
			MULT_79(2)<=signed(DIN_79_8)*signed(FMAP_3_79);
			MULT_80(2)<=signed(DIN_80_8)*signed(FMAP_3_80);
			MULT_81(2)<=signed(DIN_81_8)*signed(FMAP_3_81);
			MULT_82(2)<=signed(DIN_82_8)*signed(FMAP_3_82);
			MULT_83(2)<=signed(DIN_83_8)*signed(FMAP_3_83);
			MULT_84(2)<=signed(DIN_84_8)*signed(FMAP_3_84);

			MULT_1(3)<=signed(DIN_1_8)*signed(FMAP_4_1);
			MULT_2(3)<=signed(DIN_2_8)*signed(FMAP_4_2);
			MULT_3(3)<=signed(DIN_3_8)*signed(FMAP_4_3);
			MULT_4(3)<=signed(DIN_4_8)*signed(FMAP_4_4);
			MULT_5(3)<=signed(DIN_5_8)*signed(FMAP_4_5);
			MULT_6(3)<=signed(DIN_6_8)*signed(FMAP_4_6);
			MULT_7(3)<=signed(DIN_7_8)*signed(FMAP_4_7);
			MULT_8(3)<=signed(DIN_8_8)*signed(FMAP_4_8);
			MULT_9(3)<=signed(DIN_9_8)*signed(FMAP_4_9);
			MULT_10(3)<=signed(DIN_10_8)*signed(FMAP_4_10);
			MULT_11(3)<=signed(DIN_11_8)*signed(FMAP_4_11);
			MULT_12(3)<=signed(DIN_12_8)*signed(FMAP_4_12);
			MULT_13(3)<=signed(DIN_13_8)*signed(FMAP_4_13);
			MULT_14(3)<=signed(DIN_14_8)*signed(FMAP_4_14);
			MULT_15(3)<=signed(DIN_15_8)*signed(FMAP_4_15);
			MULT_16(3)<=signed(DIN_16_8)*signed(FMAP_4_16);
			MULT_17(3)<=signed(DIN_17_8)*signed(FMAP_4_17);
			MULT_18(3)<=signed(DIN_18_8)*signed(FMAP_4_18);
			MULT_19(3)<=signed(DIN_19_8)*signed(FMAP_4_19);
			MULT_20(3)<=signed(DIN_20_8)*signed(FMAP_4_20);
			MULT_21(3)<=signed(DIN_21_8)*signed(FMAP_4_21);
			MULT_22(3)<=signed(DIN_22_8)*signed(FMAP_4_22);
			MULT_23(3)<=signed(DIN_23_8)*signed(FMAP_4_23);
			MULT_24(3)<=signed(DIN_24_8)*signed(FMAP_4_24);
			MULT_25(3)<=signed(DIN_25_8)*signed(FMAP_4_25);
			MULT_26(3)<=signed(DIN_26_8)*signed(FMAP_4_26);
			MULT_27(3)<=signed(DIN_27_8)*signed(FMAP_4_27);
			MULT_28(3)<=signed(DIN_28_8)*signed(FMAP_4_28);
			MULT_29(3)<=signed(DIN_29_8)*signed(FMAP_4_29);
			MULT_30(3)<=signed(DIN_30_8)*signed(FMAP_4_30);
			MULT_31(3)<=signed(DIN_31_8)*signed(FMAP_4_31);
			MULT_32(3)<=signed(DIN_32_8)*signed(FMAP_4_32);
			MULT_33(3)<=signed(DIN_33_8)*signed(FMAP_4_33);
			MULT_34(3)<=signed(DIN_34_8)*signed(FMAP_4_34);
			MULT_35(3)<=signed(DIN_35_8)*signed(FMAP_4_35);
			MULT_36(3)<=signed(DIN_36_8)*signed(FMAP_4_36);
			MULT_37(3)<=signed(DIN_37_8)*signed(FMAP_4_37);
			MULT_38(3)<=signed(DIN_38_8)*signed(FMAP_4_38);
			MULT_39(3)<=signed(DIN_39_8)*signed(FMAP_4_39);
			MULT_40(3)<=signed(DIN_40_8)*signed(FMAP_4_40);
			MULT_41(3)<=signed(DIN_41_8)*signed(FMAP_4_41);
			MULT_42(3)<=signed(DIN_42_8)*signed(FMAP_4_42);
			MULT_43(3)<=signed(DIN_43_8)*signed(FMAP_4_43);
			MULT_44(3)<=signed(DIN_44_8)*signed(FMAP_4_44);
			MULT_45(3)<=signed(DIN_45_8)*signed(FMAP_4_45);
			MULT_46(3)<=signed(DIN_46_8)*signed(FMAP_4_46);
			MULT_47(3)<=signed(DIN_47_8)*signed(FMAP_4_47);
			MULT_48(3)<=signed(DIN_48_8)*signed(FMAP_4_48);
			MULT_49(3)<=signed(DIN_49_8)*signed(FMAP_4_49);
			MULT_50(3)<=signed(DIN_50_8)*signed(FMAP_4_50);
			MULT_51(3)<=signed(DIN_51_8)*signed(FMAP_4_51);
			MULT_52(3)<=signed(DIN_52_8)*signed(FMAP_4_52);
			MULT_53(3)<=signed(DIN_53_8)*signed(FMAP_4_53);
			MULT_54(3)<=signed(DIN_54_8)*signed(FMAP_4_54);
			MULT_55(3)<=signed(DIN_55_8)*signed(FMAP_4_55);
			MULT_56(3)<=signed(DIN_56_8)*signed(FMAP_4_56);
			MULT_57(3)<=signed(DIN_57_8)*signed(FMAP_4_57);
			MULT_58(3)<=signed(DIN_58_8)*signed(FMAP_4_58);
			MULT_59(3)<=signed(DIN_59_8)*signed(FMAP_4_59);
			MULT_60(3)<=signed(DIN_60_8)*signed(FMAP_4_60);
			MULT_61(3)<=signed(DIN_61_8)*signed(FMAP_4_61);
			MULT_62(3)<=signed(DIN_62_8)*signed(FMAP_4_62);
			MULT_63(3)<=signed(DIN_63_8)*signed(FMAP_4_63);
			MULT_64(3)<=signed(DIN_64_8)*signed(FMAP_4_64);
			MULT_65(3)<=signed(DIN_65_8)*signed(FMAP_4_65);
			MULT_66(3)<=signed(DIN_66_8)*signed(FMAP_4_66);
			MULT_67(3)<=signed(DIN_67_8)*signed(FMAP_4_67);
			MULT_68(3)<=signed(DIN_68_8)*signed(FMAP_4_68);
			MULT_69(3)<=signed(DIN_69_8)*signed(FMAP_4_69);
			MULT_70(3)<=signed(DIN_70_8)*signed(FMAP_4_70);
			MULT_71(3)<=signed(DIN_71_8)*signed(FMAP_4_71);
			MULT_72(3)<=signed(DIN_72_8)*signed(FMAP_4_72);
			MULT_73(3)<=signed(DIN_73_8)*signed(FMAP_4_73);
			MULT_74(3)<=signed(DIN_74_8)*signed(FMAP_4_74);
			MULT_75(3)<=signed(DIN_75_8)*signed(FMAP_4_75);
			MULT_76(3)<=signed(DIN_76_8)*signed(FMAP_4_76);
			MULT_77(3)<=signed(DIN_77_8)*signed(FMAP_4_77);
			MULT_78(3)<=signed(DIN_78_8)*signed(FMAP_4_78);
			MULT_79(3)<=signed(DIN_79_8)*signed(FMAP_4_79);
			MULT_80(3)<=signed(DIN_80_8)*signed(FMAP_4_80);
			MULT_81(3)<=signed(DIN_81_8)*signed(FMAP_4_81);
			MULT_82(3)<=signed(DIN_82_8)*signed(FMAP_4_82);
			MULT_83(3)<=signed(DIN_83_8)*signed(FMAP_4_83);
			MULT_84(3)<=signed(DIN_84_8)*signed(FMAP_4_84);

			MULT_1(4)<=signed(DIN_1_8)*signed(FMAP_5_1);
			MULT_2(4)<=signed(DIN_2_8)*signed(FMAP_5_2);
			MULT_3(4)<=signed(DIN_3_8)*signed(FMAP_5_3);
			MULT_4(4)<=signed(DIN_4_8)*signed(FMAP_5_4);
			MULT_5(4)<=signed(DIN_5_8)*signed(FMAP_5_5);
			MULT_6(4)<=signed(DIN_6_8)*signed(FMAP_5_6);
			MULT_7(4)<=signed(DIN_7_8)*signed(FMAP_5_7);
			MULT_8(4)<=signed(DIN_8_8)*signed(FMAP_5_8);
			MULT_9(4)<=signed(DIN_9_8)*signed(FMAP_5_9);
			MULT_10(4)<=signed(DIN_10_8)*signed(FMAP_5_10);
			MULT_11(4)<=signed(DIN_11_8)*signed(FMAP_5_11);
			MULT_12(4)<=signed(DIN_12_8)*signed(FMAP_5_12);
			MULT_13(4)<=signed(DIN_13_8)*signed(FMAP_5_13);
			MULT_14(4)<=signed(DIN_14_8)*signed(FMAP_5_14);
			MULT_15(4)<=signed(DIN_15_8)*signed(FMAP_5_15);
			MULT_16(4)<=signed(DIN_16_8)*signed(FMAP_5_16);
			MULT_17(4)<=signed(DIN_17_8)*signed(FMAP_5_17);
			MULT_18(4)<=signed(DIN_18_8)*signed(FMAP_5_18);
			MULT_19(4)<=signed(DIN_19_8)*signed(FMAP_5_19);
			MULT_20(4)<=signed(DIN_20_8)*signed(FMAP_5_20);
			MULT_21(4)<=signed(DIN_21_8)*signed(FMAP_5_21);
			MULT_22(4)<=signed(DIN_22_8)*signed(FMAP_5_22);
			MULT_23(4)<=signed(DIN_23_8)*signed(FMAP_5_23);
			MULT_24(4)<=signed(DIN_24_8)*signed(FMAP_5_24);
			MULT_25(4)<=signed(DIN_25_8)*signed(FMAP_5_25);
			MULT_26(4)<=signed(DIN_26_8)*signed(FMAP_5_26);
			MULT_27(4)<=signed(DIN_27_8)*signed(FMAP_5_27);
			MULT_28(4)<=signed(DIN_28_8)*signed(FMAP_5_28);
			MULT_29(4)<=signed(DIN_29_8)*signed(FMAP_5_29);
			MULT_30(4)<=signed(DIN_30_8)*signed(FMAP_5_30);
			MULT_31(4)<=signed(DIN_31_8)*signed(FMAP_5_31);
			MULT_32(4)<=signed(DIN_32_8)*signed(FMAP_5_32);
			MULT_33(4)<=signed(DIN_33_8)*signed(FMAP_5_33);
			MULT_34(4)<=signed(DIN_34_8)*signed(FMAP_5_34);
			MULT_35(4)<=signed(DIN_35_8)*signed(FMAP_5_35);
			MULT_36(4)<=signed(DIN_36_8)*signed(FMAP_5_36);
			MULT_37(4)<=signed(DIN_37_8)*signed(FMAP_5_37);
			MULT_38(4)<=signed(DIN_38_8)*signed(FMAP_5_38);
			MULT_39(4)<=signed(DIN_39_8)*signed(FMAP_5_39);
			MULT_40(4)<=signed(DIN_40_8)*signed(FMAP_5_40);
			MULT_41(4)<=signed(DIN_41_8)*signed(FMAP_5_41);
			MULT_42(4)<=signed(DIN_42_8)*signed(FMAP_5_42);
			MULT_43(4)<=signed(DIN_43_8)*signed(FMAP_5_43);
			MULT_44(4)<=signed(DIN_44_8)*signed(FMAP_5_44);
			MULT_45(4)<=signed(DIN_45_8)*signed(FMAP_5_45);
			MULT_46(4)<=signed(DIN_46_8)*signed(FMAP_5_46);
			MULT_47(4)<=signed(DIN_47_8)*signed(FMAP_5_47);
			MULT_48(4)<=signed(DIN_48_8)*signed(FMAP_5_48);
			MULT_49(4)<=signed(DIN_49_8)*signed(FMAP_5_49);
			MULT_50(4)<=signed(DIN_50_8)*signed(FMAP_5_50);
			MULT_51(4)<=signed(DIN_51_8)*signed(FMAP_5_51);
			MULT_52(4)<=signed(DIN_52_8)*signed(FMAP_5_52);
			MULT_53(4)<=signed(DIN_53_8)*signed(FMAP_5_53);
			MULT_54(4)<=signed(DIN_54_8)*signed(FMAP_5_54);
			MULT_55(4)<=signed(DIN_55_8)*signed(FMAP_5_55);
			MULT_56(4)<=signed(DIN_56_8)*signed(FMAP_5_56);
			MULT_57(4)<=signed(DIN_57_8)*signed(FMAP_5_57);
			MULT_58(4)<=signed(DIN_58_8)*signed(FMAP_5_58);
			MULT_59(4)<=signed(DIN_59_8)*signed(FMAP_5_59);
			MULT_60(4)<=signed(DIN_60_8)*signed(FMAP_5_60);
			MULT_61(4)<=signed(DIN_61_8)*signed(FMAP_5_61);
			MULT_62(4)<=signed(DIN_62_8)*signed(FMAP_5_62);
			MULT_63(4)<=signed(DIN_63_8)*signed(FMAP_5_63);
			MULT_64(4)<=signed(DIN_64_8)*signed(FMAP_5_64);
			MULT_65(4)<=signed(DIN_65_8)*signed(FMAP_5_65);
			MULT_66(4)<=signed(DIN_66_8)*signed(FMAP_5_66);
			MULT_67(4)<=signed(DIN_67_8)*signed(FMAP_5_67);
			MULT_68(4)<=signed(DIN_68_8)*signed(FMAP_5_68);
			MULT_69(4)<=signed(DIN_69_8)*signed(FMAP_5_69);
			MULT_70(4)<=signed(DIN_70_8)*signed(FMAP_5_70);
			MULT_71(4)<=signed(DIN_71_8)*signed(FMAP_5_71);
			MULT_72(4)<=signed(DIN_72_8)*signed(FMAP_5_72);
			MULT_73(4)<=signed(DIN_73_8)*signed(FMAP_5_73);
			MULT_74(4)<=signed(DIN_74_8)*signed(FMAP_5_74);
			MULT_75(4)<=signed(DIN_75_8)*signed(FMAP_5_75);
			MULT_76(4)<=signed(DIN_76_8)*signed(FMAP_5_76);
			MULT_77(4)<=signed(DIN_77_8)*signed(FMAP_5_77);
			MULT_78(4)<=signed(DIN_78_8)*signed(FMAP_5_78);
			MULT_79(4)<=signed(DIN_79_8)*signed(FMAP_5_79);
			MULT_80(4)<=signed(DIN_80_8)*signed(FMAP_5_80);
			MULT_81(4)<=signed(DIN_81_8)*signed(FMAP_5_81);
			MULT_82(4)<=signed(DIN_82_8)*signed(FMAP_5_82);
			MULT_83(4)<=signed(DIN_83_8)*signed(FMAP_5_83);
			MULT_84(4)<=signed(DIN_84_8)*signed(FMAP_5_84);

			MULT_1(5)<=signed(DIN_1_8)*signed(FMAP_6_1);
			MULT_2(5)<=signed(DIN_2_8)*signed(FMAP_6_2);
			MULT_3(5)<=signed(DIN_3_8)*signed(FMAP_6_3);
			MULT_4(5)<=signed(DIN_4_8)*signed(FMAP_6_4);
			MULT_5(5)<=signed(DIN_5_8)*signed(FMAP_6_5);
			MULT_6(5)<=signed(DIN_6_8)*signed(FMAP_6_6);
			MULT_7(5)<=signed(DIN_7_8)*signed(FMAP_6_7);
			MULT_8(5)<=signed(DIN_8_8)*signed(FMAP_6_8);
			MULT_9(5)<=signed(DIN_9_8)*signed(FMAP_6_9);
			MULT_10(5)<=signed(DIN_10_8)*signed(FMAP_6_10);
			MULT_11(5)<=signed(DIN_11_8)*signed(FMAP_6_11);
			MULT_12(5)<=signed(DIN_12_8)*signed(FMAP_6_12);
			MULT_13(5)<=signed(DIN_13_8)*signed(FMAP_6_13);
			MULT_14(5)<=signed(DIN_14_8)*signed(FMAP_6_14);
			MULT_15(5)<=signed(DIN_15_8)*signed(FMAP_6_15);
			MULT_16(5)<=signed(DIN_16_8)*signed(FMAP_6_16);
			MULT_17(5)<=signed(DIN_17_8)*signed(FMAP_6_17);
			MULT_18(5)<=signed(DIN_18_8)*signed(FMAP_6_18);
			MULT_19(5)<=signed(DIN_19_8)*signed(FMAP_6_19);
			MULT_20(5)<=signed(DIN_20_8)*signed(FMAP_6_20);
			MULT_21(5)<=signed(DIN_21_8)*signed(FMAP_6_21);
			MULT_22(5)<=signed(DIN_22_8)*signed(FMAP_6_22);
			MULT_23(5)<=signed(DIN_23_8)*signed(FMAP_6_23);
			MULT_24(5)<=signed(DIN_24_8)*signed(FMAP_6_24);
			MULT_25(5)<=signed(DIN_25_8)*signed(FMAP_6_25);
			MULT_26(5)<=signed(DIN_26_8)*signed(FMAP_6_26);
			MULT_27(5)<=signed(DIN_27_8)*signed(FMAP_6_27);
			MULT_28(5)<=signed(DIN_28_8)*signed(FMAP_6_28);
			MULT_29(5)<=signed(DIN_29_8)*signed(FMAP_6_29);
			MULT_30(5)<=signed(DIN_30_8)*signed(FMAP_6_30);
			MULT_31(5)<=signed(DIN_31_8)*signed(FMAP_6_31);
			MULT_32(5)<=signed(DIN_32_8)*signed(FMAP_6_32);
			MULT_33(5)<=signed(DIN_33_8)*signed(FMAP_6_33);
			MULT_34(5)<=signed(DIN_34_8)*signed(FMAP_6_34);
			MULT_35(5)<=signed(DIN_35_8)*signed(FMAP_6_35);
			MULT_36(5)<=signed(DIN_36_8)*signed(FMAP_6_36);
			MULT_37(5)<=signed(DIN_37_8)*signed(FMAP_6_37);
			MULT_38(5)<=signed(DIN_38_8)*signed(FMAP_6_38);
			MULT_39(5)<=signed(DIN_39_8)*signed(FMAP_6_39);
			MULT_40(5)<=signed(DIN_40_8)*signed(FMAP_6_40);
			MULT_41(5)<=signed(DIN_41_8)*signed(FMAP_6_41);
			MULT_42(5)<=signed(DIN_42_8)*signed(FMAP_6_42);
			MULT_43(5)<=signed(DIN_43_8)*signed(FMAP_6_43);
			MULT_44(5)<=signed(DIN_44_8)*signed(FMAP_6_44);
			MULT_45(5)<=signed(DIN_45_8)*signed(FMAP_6_45);
			MULT_46(5)<=signed(DIN_46_8)*signed(FMAP_6_46);
			MULT_47(5)<=signed(DIN_47_8)*signed(FMAP_6_47);
			MULT_48(5)<=signed(DIN_48_8)*signed(FMAP_6_48);
			MULT_49(5)<=signed(DIN_49_8)*signed(FMAP_6_49);
			MULT_50(5)<=signed(DIN_50_8)*signed(FMAP_6_50);
			MULT_51(5)<=signed(DIN_51_8)*signed(FMAP_6_51);
			MULT_52(5)<=signed(DIN_52_8)*signed(FMAP_6_52);
			MULT_53(5)<=signed(DIN_53_8)*signed(FMAP_6_53);
			MULT_54(5)<=signed(DIN_54_8)*signed(FMAP_6_54);
			MULT_55(5)<=signed(DIN_55_8)*signed(FMAP_6_55);
			MULT_56(5)<=signed(DIN_56_8)*signed(FMAP_6_56);
			MULT_57(5)<=signed(DIN_57_8)*signed(FMAP_6_57);
			MULT_58(5)<=signed(DIN_58_8)*signed(FMAP_6_58);
			MULT_59(5)<=signed(DIN_59_8)*signed(FMAP_6_59);
			MULT_60(5)<=signed(DIN_60_8)*signed(FMAP_6_60);
			MULT_61(5)<=signed(DIN_61_8)*signed(FMAP_6_61);
			MULT_62(5)<=signed(DIN_62_8)*signed(FMAP_6_62);
			MULT_63(5)<=signed(DIN_63_8)*signed(FMAP_6_63);
			MULT_64(5)<=signed(DIN_64_8)*signed(FMAP_6_64);
			MULT_65(5)<=signed(DIN_65_8)*signed(FMAP_6_65);
			MULT_66(5)<=signed(DIN_66_8)*signed(FMAP_6_66);
			MULT_67(5)<=signed(DIN_67_8)*signed(FMAP_6_67);
			MULT_68(5)<=signed(DIN_68_8)*signed(FMAP_6_68);
			MULT_69(5)<=signed(DIN_69_8)*signed(FMAP_6_69);
			MULT_70(5)<=signed(DIN_70_8)*signed(FMAP_6_70);
			MULT_71(5)<=signed(DIN_71_8)*signed(FMAP_6_71);
			MULT_72(5)<=signed(DIN_72_8)*signed(FMAP_6_72);
			MULT_73(5)<=signed(DIN_73_8)*signed(FMAP_6_73);
			MULT_74(5)<=signed(DIN_74_8)*signed(FMAP_6_74);
			MULT_75(5)<=signed(DIN_75_8)*signed(FMAP_6_75);
			MULT_76(5)<=signed(DIN_76_8)*signed(FMAP_6_76);
			MULT_77(5)<=signed(DIN_77_8)*signed(FMAP_6_77);
			MULT_78(5)<=signed(DIN_78_8)*signed(FMAP_6_78);
			MULT_79(5)<=signed(DIN_79_8)*signed(FMAP_6_79);
			MULT_80(5)<=signed(DIN_80_8)*signed(FMAP_6_80);
			MULT_81(5)<=signed(DIN_81_8)*signed(FMAP_6_81);
			MULT_82(5)<=signed(DIN_82_8)*signed(FMAP_6_82);
			MULT_83(5)<=signed(DIN_83_8)*signed(FMAP_6_83);
			MULT_84(5)<=signed(DIN_84_8)*signed(FMAP_6_84);

			MULT_1(6)<=signed(DIN_1_8)*signed(FMAP_7_1);
			MULT_2(6)<=signed(DIN_2_8)*signed(FMAP_7_2);
			MULT_3(6)<=signed(DIN_3_8)*signed(FMAP_7_3);
			MULT_4(6)<=signed(DIN_4_8)*signed(FMAP_7_4);
			MULT_5(6)<=signed(DIN_5_8)*signed(FMAP_7_5);
			MULT_6(6)<=signed(DIN_6_8)*signed(FMAP_7_6);
			MULT_7(6)<=signed(DIN_7_8)*signed(FMAP_7_7);
			MULT_8(6)<=signed(DIN_8_8)*signed(FMAP_7_8);
			MULT_9(6)<=signed(DIN_9_8)*signed(FMAP_7_9);
			MULT_10(6)<=signed(DIN_10_8)*signed(FMAP_7_10);
			MULT_11(6)<=signed(DIN_11_8)*signed(FMAP_7_11);
			MULT_12(6)<=signed(DIN_12_8)*signed(FMAP_7_12);
			MULT_13(6)<=signed(DIN_13_8)*signed(FMAP_7_13);
			MULT_14(6)<=signed(DIN_14_8)*signed(FMAP_7_14);
			MULT_15(6)<=signed(DIN_15_8)*signed(FMAP_7_15);
			MULT_16(6)<=signed(DIN_16_8)*signed(FMAP_7_16);
			MULT_17(6)<=signed(DIN_17_8)*signed(FMAP_7_17);
			MULT_18(6)<=signed(DIN_18_8)*signed(FMAP_7_18);
			MULT_19(6)<=signed(DIN_19_8)*signed(FMAP_7_19);
			MULT_20(6)<=signed(DIN_20_8)*signed(FMAP_7_20);
			MULT_21(6)<=signed(DIN_21_8)*signed(FMAP_7_21);
			MULT_22(6)<=signed(DIN_22_8)*signed(FMAP_7_22);
			MULT_23(6)<=signed(DIN_23_8)*signed(FMAP_7_23);
			MULT_24(6)<=signed(DIN_24_8)*signed(FMAP_7_24);
			MULT_25(6)<=signed(DIN_25_8)*signed(FMAP_7_25);
			MULT_26(6)<=signed(DIN_26_8)*signed(FMAP_7_26);
			MULT_27(6)<=signed(DIN_27_8)*signed(FMAP_7_27);
			MULT_28(6)<=signed(DIN_28_8)*signed(FMAP_7_28);
			MULT_29(6)<=signed(DIN_29_8)*signed(FMAP_7_29);
			MULT_30(6)<=signed(DIN_30_8)*signed(FMAP_7_30);
			MULT_31(6)<=signed(DIN_31_8)*signed(FMAP_7_31);
			MULT_32(6)<=signed(DIN_32_8)*signed(FMAP_7_32);
			MULT_33(6)<=signed(DIN_33_8)*signed(FMAP_7_33);
			MULT_34(6)<=signed(DIN_34_8)*signed(FMAP_7_34);
			MULT_35(6)<=signed(DIN_35_8)*signed(FMAP_7_35);
			MULT_36(6)<=signed(DIN_36_8)*signed(FMAP_7_36);
			MULT_37(6)<=signed(DIN_37_8)*signed(FMAP_7_37);
			MULT_38(6)<=signed(DIN_38_8)*signed(FMAP_7_38);
			MULT_39(6)<=signed(DIN_39_8)*signed(FMAP_7_39);
			MULT_40(6)<=signed(DIN_40_8)*signed(FMAP_7_40);
			MULT_41(6)<=signed(DIN_41_8)*signed(FMAP_7_41);
			MULT_42(6)<=signed(DIN_42_8)*signed(FMAP_7_42);
			MULT_43(6)<=signed(DIN_43_8)*signed(FMAP_7_43);
			MULT_44(6)<=signed(DIN_44_8)*signed(FMAP_7_44);
			MULT_45(6)<=signed(DIN_45_8)*signed(FMAP_7_45);
			MULT_46(6)<=signed(DIN_46_8)*signed(FMAP_7_46);
			MULT_47(6)<=signed(DIN_47_8)*signed(FMAP_7_47);
			MULT_48(6)<=signed(DIN_48_8)*signed(FMAP_7_48);
			MULT_49(6)<=signed(DIN_49_8)*signed(FMAP_7_49);
			MULT_50(6)<=signed(DIN_50_8)*signed(FMAP_7_50);
			MULT_51(6)<=signed(DIN_51_8)*signed(FMAP_7_51);
			MULT_52(6)<=signed(DIN_52_8)*signed(FMAP_7_52);
			MULT_53(6)<=signed(DIN_53_8)*signed(FMAP_7_53);
			MULT_54(6)<=signed(DIN_54_8)*signed(FMAP_7_54);
			MULT_55(6)<=signed(DIN_55_8)*signed(FMAP_7_55);
			MULT_56(6)<=signed(DIN_56_8)*signed(FMAP_7_56);
			MULT_57(6)<=signed(DIN_57_8)*signed(FMAP_7_57);
			MULT_58(6)<=signed(DIN_58_8)*signed(FMAP_7_58);
			MULT_59(6)<=signed(DIN_59_8)*signed(FMAP_7_59);
			MULT_60(6)<=signed(DIN_60_8)*signed(FMAP_7_60);
			MULT_61(6)<=signed(DIN_61_8)*signed(FMAP_7_61);
			MULT_62(6)<=signed(DIN_62_8)*signed(FMAP_7_62);
			MULT_63(6)<=signed(DIN_63_8)*signed(FMAP_7_63);
			MULT_64(6)<=signed(DIN_64_8)*signed(FMAP_7_64);
			MULT_65(6)<=signed(DIN_65_8)*signed(FMAP_7_65);
			MULT_66(6)<=signed(DIN_66_8)*signed(FMAP_7_66);
			MULT_67(6)<=signed(DIN_67_8)*signed(FMAP_7_67);
			MULT_68(6)<=signed(DIN_68_8)*signed(FMAP_7_68);
			MULT_69(6)<=signed(DIN_69_8)*signed(FMAP_7_69);
			MULT_70(6)<=signed(DIN_70_8)*signed(FMAP_7_70);
			MULT_71(6)<=signed(DIN_71_8)*signed(FMAP_7_71);
			MULT_72(6)<=signed(DIN_72_8)*signed(FMAP_7_72);
			MULT_73(6)<=signed(DIN_73_8)*signed(FMAP_7_73);
			MULT_74(6)<=signed(DIN_74_8)*signed(FMAP_7_74);
			MULT_75(6)<=signed(DIN_75_8)*signed(FMAP_7_75);
			MULT_76(6)<=signed(DIN_76_8)*signed(FMAP_7_76);
			MULT_77(6)<=signed(DIN_77_8)*signed(FMAP_7_77);
			MULT_78(6)<=signed(DIN_78_8)*signed(FMAP_7_78);
			MULT_79(6)<=signed(DIN_79_8)*signed(FMAP_7_79);
			MULT_80(6)<=signed(DIN_80_8)*signed(FMAP_7_80);
			MULT_81(6)<=signed(DIN_81_8)*signed(FMAP_7_81);
			MULT_82(6)<=signed(DIN_82_8)*signed(FMAP_7_82);
			MULT_83(6)<=signed(DIN_83_8)*signed(FMAP_7_83);
			MULT_84(6)<=signed(DIN_84_8)*signed(FMAP_7_84);

			MULT_1(7)<=signed(DIN_1_8)*signed(FMAP_8_1);
			MULT_2(7)<=signed(DIN_2_8)*signed(FMAP_8_2);
			MULT_3(7)<=signed(DIN_3_8)*signed(FMAP_8_3);
			MULT_4(7)<=signed(DIN_4_8)*signed(FMAP_8_4);
			MULT_5(7)<=signed(DIN_5_8)*signed(FMAP_8_5);
			MULT_6(7)<=signed(DIN_6_8)*signed(FMAP_8_6);
			MULT_7(7)<=signed(DIN_7_8)*signed(FMAP_8_7);
			MULT_8(7)<=signed(DIN_8_8)*signed(FMAP_8_8);
			MULT_9(7)<=signed(DIN_9_8)*signed(FMAP_8_9);
			MULT_10(7)<=signed(DIN_10_8)*signed(FMAP_8_10);
			MULT_11(7)<=signed(DIN_11_8)*signed(FMAP_8_11);
			MULT_12(7)<=signed(DIN_12_8)*signed(FMAP_8_12);
			MULT_13(7)<=signed(DIN_13_8)*signed(FMAP_8_13);
			MULT_14(7)<=signed(DIN_14_8)*signed(FMAP_8_14);
			MULT_15(7)<=signed(DIN_15_8)*signed(FMAP_8_15);
			MULT_16(7)<=signed(DIN_16_8)*signed(FMAP_8_16);
			MULT_17(7)<=signed(DIN_17_8)*signed(FMAP_8_17);
			MULT_18(7)<=signed(DIN_18_8)*signed(FMAP_8_18);
			MULT_19(7)<=signed(DIN_19_8)*signed(FMAP_8_19);
			MULT_20(7)<=signed(DIN_20_8)*signed(FMAP_8_20);
			MULT_21(7)<=signed(DIN_21_8)*signed(FMAP_8_21);
			MULT_22(7)<=signed(DIN_22_8)*signed(FMAP_8_22);
			MULT_23(7)<=signed(DIN_23_8)*signed(FMAP_8_23);
			MULT_24(7)<=signed(DIN_24_8)*signed(FMAP_8_24);
			MULT_25(7)<=signed(DIN_25_8)*signed(FMAP_8_25);
			MULT_26(7)<=signed(DIN_26_8)*signed(FMAP_8_26);
			MULT_27(7)<=signed(DIN_27_8)*signed(FMAP_8_27);
			MULT_28(7)<=signed(DIN_28_8)*signed(FMAP_8_28);
			MULT_29(7)<=signed(DIN_29_8)*signed(FMAP_8_29);
			MULT_30(7)<=signed(DIN_30_8)*signed(FMAP_8_30);
			MULT_31(7)<=signed(DIN_31_8)*signed(FMAP_8_31);
			MULT_32(7)<=signed(DIN_32_8)*signed(FMAP_8_32);
			MULT_33(7)<=signed(DIN_33_8)*signed(FMAP_8_33);
			MULT_34(7)<=signed(DIN_34_8)*signed(FMAP_8_34);
			MULT_35(7)<=signed(DIN_35_8)*signed(FMAP_8_35);
			MULT_36(7)<=signed(DIN_36_8)*signed(FMAP_8_36);
			MULT_37(7)<=signed(DIN_37_8)*signed(FMAP_8_37);
			MULT_38(7)<=signed(DIN_38_8)*signed(FMAP_8_38);
			MULT_39(7)<=signed(DIN_39_8)*signed(FMAP_8_39);
			MULT_40(7)<=signed(DIN_40_8)*signed(FMAP_8_40);
			MULT_41(7)<=signed(DIN_41_8)*signed(FMAP_8_41);
			MULT_42(7)<=signed(DIN_42_8)*signed(FMAP_8_42);
			MULT_43(7)<=signed(DIN_43_8)*signed(FMAP_8_43);
			MULT_44(7)<=signed(DIN_44_8)*signed(FMAP_8_44);
			MULT_45(7)<=signed(DIN_45_8)*signed(FMAP_8_45);
			MULT_46(7)<=signed(DIN_46_8)*signed(FMAP_8_46);
			MULT_47(7)<=signed(DIN_47_8)*signed(FMAP_8_47);
			MULT_48(7)<=signed(DIN_48_8)*signed(FMAP_8_48);
			MULT_49(7)<=signed(DIN_49_8)*signed(FMAP_8_49);
			MULT_50(7)<=signed(DIN_50_8)*signed(FMAP_8_50);
			MULT_51(7)<=signed(DIN_51_8)*signed(FMAP_8_51);
			MULT_52(7)<=signed(DIN_52_8)*signed(FMAP_8_52);
			MULT_53(7)<=signed(DIN_53_8)*signed(FMAP_8_53);
			MULT_54(7)<=signed(DIN_54_8)*signed(FMAP_8_54);
			MULT_55(7)<=signed(DIN_55_8)*signed(FMAP_8_55);
			MULT_56(7)<=signed(DIN_56_8)*signed(FMAP_8_56);
			MULT_57(7)<=signed(DIN_57_8)*signed(FMAP_8_57);
			MULT_58(7)<=signed(DIN_58_8)*signed(FMAP_8_58);
			MULT_59(7)<=signed(DIN_59_8)*signed(FMAP_8_59);
			MULT_60(7)<=signed(DIN_60_8)*signed(FMAP_8_60);
			MULT_61(7)<=signed(DIN_61_8)*signed(FMAP_8_61);
			MULT_62(7)<=signed(DIN_62_8)*signed(FMAP_8_62);
			MULT_63(7)<=signed(DIN_63_8)*signed(FMAP_8_63);
			MULT_64(7)<=signed(DIN_64_8)*signed(FMAP_8_64);
			MULT_65(7)<=signed(DIN_65_8)*signed(FMAP_8_65);
			MULT_66(7)<=signed(DIN_66_8)*signed(FMAP_8_66);
			MULT_67(7)<=signed(DIN_67_8)*signed(FMAP_8_67);
			MULT_68(7)<=signed(DIN_68_8)*signed(FMAP_8_68);
			MULT_69(7)<=signed(DIN_69_8)*signed(FMAP_8_69);
			MULT_70(7)<=signed(DIN_70_8)*signed(FMAP_8_70);
			MULT_71(7)<=signed(DIN_71_8)*signed(FMAP_8_71);
			MULT_72(7)<=signed(DIN_72_8)*signed(FMAP_8_72);
			MULT_73(7)<=signed(DIN_73_8)*signed(FMAP_8_73);
			MULT_74(7)<=signed(DIN_74_8)*signed(FMAP_8_74);
			MULT_75(7)<=signed(DIN_75_8)*signed(FMAP_8_75);
			MULT_76(7)<=signed(DIN_76_8)*signed(FMAP_8_76);
			MULT_77(7)<=signed(DIN_77_8)*signed(FMAP_8_77);
			MULT_78(7)<=signed(DIN_78_8)*signed(FMAP_8_78);
			MULT_79(7)<=signed(DIN_79_8)*signed(FMAP_8_79);
			MULT_80(7)<=signed(DIN_80_8)*signed(FMAP_8_80);
			MULT_81(7)<=signed(DIN_81_8)*signed(FMAP_8_81);
			MULT_82(7)<=signed(DIN_82_8)*signed(FMAP_8_82);
			MULT_83(7)<=signed(DIN_83_8)*signed(FMAP_8_83);
			MULT_84(7)<=signed(DIN_84_8)*signed(FMAP_8_84);

			MULT_1(8)<=signed(DIN_1_8)*signed(FMAP_9_1);
			MULT_2(8)<=signed(DIN_2_8)*signed(FMAP_9_2);
			MULT_3(8)<=signed(DIN_3_8)*signed(FMAP_9_3);
			MULT_4(8)<=signed(DIN_4_8)*signed(FMAP_9_4);
			MULT_5(8)<=signed(DIN_5_8)*signed(FMAP_9_5);
			MULT_6(8)<=signed(DIN_6_8)*signed(FMAP_9_6);
			MULT_7(8)<=signed(DIN_7_8)*signed(FMAP_9_7);
			MULT_8(8)<=signed(DIN_8_8)*signed(FMAP_9_8);
			MULT_9(8)<=signed(DIN_9_8)*signed(FMAP_9_9);
			MULT_10(8)<=signed(DIN_10_8)*signed(FMAP_9_10);
			MULT_11(8)<=signed(DIN_11_8)*signed(FMAP_9_11);
			MULT_12(8)<=signed(DIN_12_8)*signed(FMAP_9_12);
			MULT_13(8)<=signed(DIN_13_8)*signed(FMAP_9_13);
			MULT_14(8)<=signed(DIN_14_8)*signed(FMAP_9_14);
			MULT_15(8)<=signed(DIN_15_8)*signed(FMAP_9_15);
			MULT_16(8)<=signed(DIN_16_8)*signed(FMAP_9_16);
			MULT_17(8)<=signed(DIN_17_8)*signed(FMAP_9_17);
			MULT_18(8)<=signed(DIN_18_8)*signed(FMAP_9_18);
			MULT_19(8)<=signed(DIN_19_8)*signed(FMAP_9_19);
			MULT_20(8)<=signed(DIN_20_8)*signed(FMAP_9_20);
			MULT_21(8)<=signed(DIN_21_8)*signed(FMAP_9_21);
			MULT_22(8)<=signed(DIN_22_8)*signed(FMAP_9_22);
			MULT_23(8)<=signed(DIN_23_8)*signed(FMAP_9_23);
			MULT_24(8)<=signed(DIN_24_8)*signed(FMAP_9_24);
			MULT_25(8)<=signed(DIN_25_8)*signed(FMAP_9_25);
			MULT_26(8)<=signed(DIN_26_8)*signed(FMAP_9_26);
			MULT_27(8)<=signed(DIN_27_8)*signed(FMAP_9_27);
			MULT_28(8)<=signed(DIN_28_8)*signed(FMAP_9_28);
			MULT_29(8)<=signed(DIN_29_8)*signed(FMAP_9_29);
			MULT_30(8)<=signed(DIN_30_8)*signed(FMAP_9_30);
			MULT_31(8)<=signed(DIN_31_8)*signed(FMAP_9_31);
			MULT_32(8)<=signed(DIN_32_8)*signed(FMAP_9_32);
			MULT_33(8)<=signed(DIN_33_8)*signed(FMAP_9_33);
			MULT_34(8)<=signed(DIN_34_8)*signed(FMAP_9_34);
			MULT_35(8)<=signed(DIN_35_8)*signed(FMAP_9_35);
			MULT_36(8)<=signed(DIN_36_8)*signed(FMAP_9_36);
			MULT_37(8)<=signed(DIN_37_8)*signed(FMAP_9_37);
			MULT_38(8)<=signed(DIN_38_8)*signed(FMAP_9_38);
			MULT_39(8)<=signed(DIN_39_8)*signed(FMAP_9_39);
			MULT_40(8)<=signed(DIN_40_8)*signed(FMAP_9_40);
			MULT_41(8)<=signed(DIN_41_8)*signed(FMAP_9_41);
			MULT_42(8)<=signed(DIN_42_8)*signed(FMAP_9_42);
			MULT_43(8)<=signed(DIN_43_8)*signed(FMAP_9_43);
			MULT_44(8)<=signed(DIN_44_8)*signed(FMAP_9_44);
			MULT_45(8)<=signed(DIN_45_8)*signed(FMAP_9_45);
			MULT_46(8)<=signed(DIN_46_8)*signed(FMAP_9_46);
			MULT_47(8)<=signed(DIN_47_8)*signed(FMAP_9_47);
			MULT_48(8)<=signed(DIN_48_8)*signed(FMAP_9_48);
			MULT_49(8)<=signed(DIN_49_8)*signed(FMAP_9_49);
			MULT_50(8)<=signed(DIN_50_8)*signed(FMAP_9_50);
			MULT_51(8)<=signed(DIN_51_8)*signed(FMAP_9_51);
			MULT_52(8)<=signed(DIN_52_8)*signed(FMAP_9_52);
			MULT_53(8)<=signed(DIN_53_8)*signed(FMAP_9_53);
			MULT_54(8)<=signed(DIN_54_8)*signed(FMAP_9_54);
			MULT_55(8)<=signed(DIN_55_8)*signed(FMAP_9_55);
			MULT_56(8)<=signed(DIN_56_8)*signed(FMAP_9_56);
			MULT_57(8)<=signed(DIN_57_8)*signed(FMAP_9_57);
			MULT_58(8)<=signed(DIN_58_8)*signed(FMAP_9_58);
			MULT_59(8)<=signed(DIN_59_8)*signed(FMAP_9_59);
			MULT_60(8)<=signed(DIN_60_8)*signed(FMAP_9_60);
			MULT_61(8)<=signed(DIN_61_8)*signed(FMAP_9_61);
			MULT_62(8)<=signed(DIN_62_8)*signed(FMAP_9_62);
			MULT_63(8)<=signed(DIN_63_8)*signed(FMAP_9_63);
			MULT_64(8)<=signed(DIN_64_8)*signed(FMAP_9_64);
			MULT_65(8)<=signed(DIN_65_8)*signed(FMAP_9_65);
			MULT_66(8)<=signed(DIN_66_8)*signed(FMAP_9_66);
			MULT_67(8)<=signed(DIN_67_8)*signed(FMAP_9_67);
			MULT_68(8)<=signed(DIN_68_8)*signed(FMAP_9_68);
			MULT_69(8)<=signed(DIN_69_8)*signed(FMAP_9_69);
			MULT_70(8)<=signed(DIN_70_8)*signed(FMAP_9_70);
			MULT_71(8)<=signed(DIN_71_8)*signed(FMAP_9_71);
			MULT_72(8)<=signed(DIN_72_8)*signed(FMAP_9_72);
			MULT_73(8)<=signed(DIN_73_8)*signed(FMAP_9_73);
			MULT_74(8)<=signed(DIN_74_8)*signed(FMAP_9_74);
			MULT_75(8)<=signed(DIN_75_8)*signed(FMAP_9_75);
			MULT_76(8)<=signed(DIN_76_8)*signed(FMAP_9_76);
			MULT_77(8)<=signed(DIN_77_8)*signed(FMAP_9_77);
			MULT_78(8)<=signed(DIN_78_8)*signed(FMAP_9_78);
			MULT_79(8)<=signed(DIN_79_8)*signed(FMAP_9_79);
			MULT_80(8)<=signed(DIN_80_8)*signed(FMAP_9_80);
			MULT_81(8)<=signed(DIN_81_8)*signed(FMAP_9_81);
			MULT_82(8)<=signed(DIN_82_8)*signed(FMAP_9_82);
			MULT_83(8)<=signed(DIN_83_8)*signed(FMAP_9_83);
			MULT_84(8)<=signed(DIN_84_8)*signed(FMAP_9_84);

			MULT_1(9)<=signed(DIN_1_8)*signed(FMAP_10_1);
			MULT_2(9)<=signed(DIN_2_8)*signed(FMAP_10_2);
			MULT_3(9)<=signed(DIN_3_8)*signed(FMAP_10_3);
			MULT_4(9)<=signed(DIN_4_8)*signed(FMAP_10_4);
			MULT_5(9)<=signed(DIN_5_8)*signed(FMAP_10_5);
			MULT_6(9)<=signed(DIN_6_8)*signed(FMAP_10_6);
			MULT_7(9)<=signed(DIN_7_8)*signed(FMAP_10_7);
			MULT_8(9)<=signed(DIN_8_8)*signed(FMAP_10_8);
			MULT_9(9)<=signed(DIN_9_8)*signed(FMAP_10_9);
			MULT_10(9)<=signed(DIN_10_8)*signed(FMAP_10_10);
			MULT_11(9)<=signed(DIN_11_8)*signed(FMAP_10_11);
			MULT_12(9)<=signed(DIN_12_8)*signed(FMAP_10_12);
			MULT_13(9)<=signed(DIN_13_8)*signed(FMAP_10_13);
			MULT_14(9)<=signed(DIN_14_8)*signed(FMAP_10_14);
			MULT_15(9)<=signed(DIN_15_8)*signed(FMAP_10_15);
			MULT_16(9)<=signed(DIN_16_8)*signed(FMAP_10_16);
			MULT_17(9)<=signed(DIN_17_8)*signed(FMAP_10_17);
			MULT_18(9)<=signed(DIN_18_8)*signed(FMAP_10_18);
			MULT_19(9)<=signed(DIN_19_8)*signed(FMAP_10_19);
			MULT_20(9)<=signed(DIN_20_8)*signed(FMAP_10_20);
			MULT_21(9)<=signed(DIN_21_8)*signed(FMAP_10_21);
			MULT_22(9)<=signed(DIN_22_8)*signed(FMAP_10_22);
			MULT_23(9)<=signed(DIN_23_8)*signed(FMAP_10_23);
			MULT_24(9)<=signed(DIN_24_8)*signed(FMAP_10_24);
			MULT_25(9)<=signed(DIN_25_8)*signed(FMAP_10_25);
			MULT_26(9)<=signed(DIN_26_8)*signed(FMAP_10_26);
			MULT_27(9)<=signed(DIN_27_8)*signed(FMAP_10_27);
			MULT_28(9)<=signed(DIN_28_8)*signed(FMAP_10_28);
			MULT_29(9)<=signed(DIN_29_8)*signed(FMAP_10_29);
			MULT_30(9)<=signed(DIN_30_8)*signed(FMAP_10_30);
			MULT_31(9)<=signed(DIN_31_8)*signed(FMAP_10_31);
			MULT_32(9)<=signed(DIN_32_8)*signed(FMAP_10_32);
			MULT_33(9)<=signed(DIN_33_8)*signed(FMAP_10_33);
			MULT_34(9)<=signed(DIN_34_8)*signed(FMAP_10_34);
			MULT_35(9)<=signed(DIN_35_8)*signed(FMAP_10_35);
			MULT_36(9)<=signed(DIN_36_8)*signed(FMAP_10_36);
			MULT_37(9)<=signed(DIN_37_8)*signed(FMAP_10_37);
			MULT_38(9)<=signed(DIN_38_8)*signed(FMAP_10_38);
			MULT_39(9)<=signed(DIN_39_8)*signed(FMAP_10_39);
			MULT_40(9)<=signed(DIN_40_8)*signed(FMAP_10_40);
			MULT_41(9)<=signed(DIN_41_8)*signed(FMAP_10_41);
			MULT_42(9)<=signed(DIN_42_8)*signed(FMAP_10_42);
			MULT_43(9)<=signed(DIN_43_8)*signed(FMAP_10_43);
			MULT_44(9)<=signed(DIN_44_8)*signed(FMAP_10_44);
			MULT_45(9)<=signed(DIN_45_8)*signed(FMAP_10_45);
			MULT_46(9)<=signed(DIN_46_8)*signed(FMAP_10_46);
			MULT_47(9)<=signed(DIN_47_8)*signed(FMAP_10_47);
			MULT_48(9)<=signed(DIN_48_8)*signed(FMAP_10_48);
			MULT_49(9)<=signed(DIN_49_8)*signed(FMAP_10_49);
			MULT_50(9)<=signed(DIN_50_8)*signed(FMAP_10_50);
			MULT_51(9)<=signed(DIN_51_8)*signed(FMAP_10_51);
			MULT_52(9)<=signed(DIN_52_8)*signed(FMAP_10_52);
			MULT_53(9)<=signed(DIN_53_8)*signed(FMAP_10_53);
			MULT_54(9)<=signed(DIN_54_8)*signed(FMAP_10_54);
			MULT_55(9)<=signed(DIN_55_8)*signed(FMAP_10_55);
			MULT_56(9)<=signed(DIN_56_8)*signed(FMAP_10_56);
			MULT_57(9)<=signed(DIN_57_8)*signed(FMAP_10_57);
			MULT_58(9)<=signed(DIN_58_8)*signed(FMAP_10_58);
			MULT_59(9)<=signed(DIN_59_8)*signed(FMAP_10_59);
			MULT_60(9)<=signed(DIN_60_8)*signed(FMAP_10_60);
			MULT_61(9)<=signed(DIN_61_8)*signed(FMAP_10_61);
			MULT_62(9)<=signed(DIN_62_8)*signed(FMAP_10_62);
			MULT_63(9)<=signed(DIN_63_8)*signed(FMAP_10_63);
			MULT_64(9)<=signed(DIN_64_8)*signed(FMAP_10_64);
			MULT_65(9)<=signed(DIN_65_8)*signed(FMAP_10_65);
			MULT_66(9)<=signed(DIN_66_8)*signed(FMAP_10_66);
			MULT_67(9)<=signed(DIN_67_8)*signed(FMAP_10_67);
			MULT_68(9)<=signed(DIN_68_8)*signed(FMAP_10_68);
			MULT_69(9)<=signed(DIN_69_8)*signed(FMAP_10_69);
			MULT_70(9)<=signed(DIN_70_8)*signed(FMAP_10_70);
			MULT_71(9)<=signed(DIN_71_8)*signed(FMAP_10_71);
			MULT_72(9)<=signed(DIN_72_8)*signed(FMAP_10_72);
			MULT_73(9)<=signed(DIN_73_8)*signed(FMAP_10_73);
			MULT_74(9)<=signed(DIN_74_8)*signed(FMAP_10_74);
			MULT_75(9)<=signed(DIN_75_8)*signed(FMAP_10_75);
			MULT_76(9)<=signed(DIN_76_8)*signed(FMAP_10_76);
			MULT_77(9)<=signed(DIN_77_8)*signed(FMAP_10_77);
			MULT_78(9)<=signed(DIN_78_8)*signed(FMAP_10_78);
			MULT_79(9)<=signed(DIN_79_8)*signed(FMAP_10_79);
			MULT_80(9)<=signed(DIN_80_8)*signed(FMAP_10_80);
			MULT_81(9)<=signed(DIN_81_8)*signed(FMAP_10_81);
			MULT_82(9)<=signed(DIN_82_8)*signed(FMAP_10_82);
			MULT_83(9)<=signed(DIN_83_8)*signed(FMAP_10_83);
			MULT_84(9)<=signed(DIN_84_8)*signed(FMAP_10_84);


                        EN_SUM_MULT_1<='1';

      -------------------------------------------- Enable MULT START --------------------------------------------				


		if EN_SUM_MULT_1 = '1' then
			------------------------------------STAGE-1--------------------------------------
			MULTS_1_1(0)<=signed(MULT_1(0)(MULT_SIZE-1) & MULT_1(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(0)(MULT_SIZE-1) & MULT_2(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(1)<=signed(MULT_1(1)(MULT_SIZE-1) & MULT_1(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(1)(MULT_SIZE-1) & MULT_2(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(2)<=signed(MULT_1(2)(MULT_SIZE-1) & MULT_1(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(2)(MULT_SIZE-1) & MULT_2(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(3)<=signed(MULT_1(3)(MULT_SIZE-1) & MULT_1(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(3)(MULT_SIZE-1) & MULT_2(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(4)<=signed(MULT_1(4)(MULT_SIZE-1) & MULT_1(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(4)(MULT_SIZE-1) & MULT_2(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(5)<=signed(MULT_1(5)(MULT_SIZE-1) & MULT_1(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(5)(MULT_SIZE-1) & MULT_2(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(6)<=signed(MULT_1(6)(MULT_SIZE-1) & MULT_1(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(6)(MULT_SIZE-1) & MULT_2(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(7)<=signed(MULT_1(7)(MULT_SIZE-1) & MULT_1(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(7)(MULT_SIZE-1) & MULT_2(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(8)<=signed(MULT_1(8)(MULT_SIZE-1) & MULT_1(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(8)(MULT_SIZE-1) & MULT_2(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(9)<=signed(MULT_1(9)(MULT_SIZE-1) & MULT_1(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(9)(MULT_SIZE-1) & MULT_2(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_2(0)<=signed(MULT_3(0)(MULT_SIZE-1) & MULT_3(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(0)(MULT_SIZE-1) & MULT_4(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(1)<=signed(MULT_3(1)(MULT_SIZE-1) & MULT_3(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(1)(MULT_SIZE-1) & MULT_4(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(2)<=signed(MULT_3(2)(MULT_SIZE-1) & MULT_3(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(2)(MULT_SIZE-1) & MULT_4(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(3)<=signed(MULT_3(3)(MULT_SIZE-1) & MULT_3(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(3)(MULT_SIZE-1) & MULT_4(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(4)<=signed(MULT_3(4)(MULT_SIZE-1) & MULT_3(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(4)(MULT_SIZE-1) & MULT_4(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(5)<=signed(MULT_3(5)(MULT_SIZE-1) & MULT_3(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(5)(MULT_SIZE-1) & MULT_4(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(6)<=signed(MULT_3(6)(MULT_SIZE-1) & MULT_3(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(6)(MULT_SIZE-1) & MULT_4(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(7)<=signed(MULT_3(7)(MULT_SIZE-1) & MULT_3(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(7)(MULT_SIZE-1) & MULT_4(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(8)<=signed(MULT_3(8)(MULT_SIZE-1) & MULT_3(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(8)(MULT_SIZE-1) & MULT_4(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(9)<=signed(MULT_3(9)(MULT_SIZE-1) & MULT_3(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(9)(MULT_SIZE-1) & MULT_4(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_3(0)<=signed(MULT_5(0)(MULT_SIZE-1) & MULT_5(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(0)(MULT_SIZE-1) & MULT_6(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(1)<=signed(MULT_5(1)(MULT_SIZE-1) & MULT_5(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(1)(MULT_SIZE-1) & MULT_6(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(2)<=signed(MULT_5(2)(MULT_SIZE-1) & MULT_5(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(2)(MULT_SIZE-1) & MULT_6(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(3)<=signed(MULT_5(3)(MULT_SIZE-1) & MULT_5(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(3)(MULT_SIZE-1) & MULT_6(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(4)<=signed(MULT_5(4)(MULT_SIZE-1) & MULT_5(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(4)(MULT_SIZE-1) & MULT_6(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(5)<=signed(MULT_5(5)(MULT_SIZE-1) & MULT_5(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(5)(MULT_SIZE-1) & MULT_6(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(6)<=signed(MULT_5(6)(MULT_SIZE-1) & MULT_5(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(6)(MULT_SIZE-1) & MULT_6(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(7)<=signed(MULT_5(7)(MULT_SIZE-1) & MULT_5(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(7)(MULT_SIZE-1) & MULT_6(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(8)<=signed(MULT_5(8)(MULT_SIZE-1) & MULT_5(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(8)(MULT_SIZE-1) & MULT_6(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(9)<=signed(MULT_5(9)(MULT_SIZE-1) & MULT_5(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(9)(MULT_SIZE-1) & MULT_6(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_4(0)<=signed(MULT_7(0)(MULT_SIZE-1) & MULT_7(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(0)(MULT_SIZE-1) & MULT_8(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(1)<=signed(MULT_7(1)(MULT_SIZE-1) & MULT_7(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(1)(MULT_SIZE-1) & MULT_8(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(2)<=signed(MULT_7(2)(MULT_SIZE-1) & MULT_7(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(2)(MULT_SIZE-1) & MULT_8(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(3)<=signed(MULT_7(3)(MULT_SIZE-1) & MULT_7(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(3)(MULT_SIZE-1) & MULT_8(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(4)<=signed(MULT_7(4)(MULT_SIZE-1) & MULT_7(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(4)(MULT_SIZE-1) & MULT_8(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(5)<=signed(MULT_7(5)(MULT_SIZE-1) & MULT_7(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(5)(MULT_SIZE-1) & MULT_8(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(6)<=signed(MULT_7(6)(MULT_SIZE-1) & MULT_7(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(6)(MULT_SIZE-1) & MULT_8(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(7)<=signed(MULT_7(7)(MULT_SIZE-1) & MULT_7(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(7)(MULT_SIZE-1) & MULT_8(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(8)<=signed(MULT_7(8)(MULT_SIZE-1) & MULT_7(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(8)(MULT_SIZE-1) & MULT_8(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(9)<=signed(MULT_7(9)(MULT_SIZE-1) & MULT_7(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(9)(MULT_SIZE-1) & MULT_8(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_5(0)<=signed(MULT_9(0)(MULT_SIZE-1) & MULT_9(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(0)(MULT_SIZE-1) & MULT_10(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(1)<=signed(MULT_9(1)(MULT_SIZE-1) & MULT_9(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(1)(MULT_SIZE-1) & MULT_10(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(2)<=signed(MULT_9(2)(MULT_SIZE-1) & MULT_9(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(2)(MULT_SIZE-1) & MULT_10(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(3)<=signed(MULT_9(3)(MULT_SIZE-1) & MULT_9(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(3)(MULT_SIZE-1) & MULT_10(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(4)<=signed(MULT_9(4)(MULT_SIZE-1) & MULT_9(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(4)(MULT_SIZE-1) & MULT_10(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(5)<=signed(MULT_9(5)(MULT_SIZE-1) & MULT_9(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(5)(MULT_SIZE-1) & MULT_10(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(6)<=signed(MULT_9(6)(MULT_SIZE-1) & MULT_9(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(6)(MULT_SIZE-1) & MULT_10(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(7)<=signed(MULT_9(7)(MULT_SIZE-1) & MULT_9(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(7)(MULT_SIZE-1) & MULT_10(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(8)<=signed(MULT_9(8)(MULT_SIZE-1) & MULT_9(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(8)(MULT_SIZE-1) & MULT_10(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(9)<=signed(MULT_9(9)(MULT_SIZE-1) & MULT_9(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(9)(MULT_SIZE-1) & MULT_10(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_6(0)<=signed(MULT_11(0)(MULT_SIZE-1) & MULT_11(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(0)(MULT_SIZE-1) & MULT_12(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(1)<=signed(MULT_11(1)(MULT_SIZE-1) & MULT_11(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(1)(MULT_SIZE-1) & MULT_12(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(2)<=signed(MULT_11(2)(MULT_SIZE-1) & MULT_11(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(2)(MULT_SIZE-1) & MULT_12(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(3)<=signed(MULT_11(3)(MULT_SIZE-1) & MULT_11(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(3)(MULT_SIZE-1) & MULT_12(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(4)<=signed(MULT_11(4)(MULT_SIZE-1) & MULT_11(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(4)(MULT_SIZE-1) & MULT_12(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(5)<=signed(MULT_11(5)(MULT_SIZE-1) & MULT_11(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(5)(MULT_SIZE-1) & MULT_12(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(6)<=signed(MULT_11(6)(MULT_SIZE-1) & MULT_11(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(6)(MULT_SIZE-1) & MULT_12(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(7)<=signed(MULT_11(7)(MULT_SIZE-1) & MULT_11(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(7)(MULT_SIZE-1) & MULT_12(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(8)<=signed(MULT_11(8)(MULT_SIZE-1) & MULT_11(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(8)(MULT_SIZE-1) & MULT_12(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(9)<=signed(MULT_11(9)(MULT_SIZE-1) & MULT_11(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(9)(MULT_SIZE-1) & MULT_12(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_7(0)<=signed(MULT_13(0)(MULT_SIZE-1) & MULT_13(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(0)(MULT_SIZE-1) & MULT_14(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(1)<=signed(MULT_13(1)(MULT_SIZE-1) & MULT_13(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(1)(MULT_SIZE-1) & MULT_14(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(2)<=signed(MULT_13(2)(MULT_SIZE-1) & MULT_13(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(2)(MULT_SIZE-1) & MULT_14(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(3)<=signed(MULT_13(3)(MULT_SIZE-1) & MULT_13(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(3)(MULT_SIZE-1) & MULT_14(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(4)<=signed(MULT_13(4)(MULT_SIZE-1) & MULT_13(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(4)(MULT_SIZE-1) & MULT_14(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(5)<=signed(MULT_13(5)(MULT_SIZE-1) & MULT_13(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(5)(MULT_SIZE-1) & MULT_14(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(6)<=signed(MULT_13(6)(MULT_SIZE-1) & MULT_13(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(6)(MULT_SIZE-1) & MULT_14(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(7)<=signed(MULT_13(7)(MULT_SIZE-1) & MULT_13(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(7)(MULT_SIZE-1) & MULT_14(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(8)<=signed(MULT_13(8)(MULT_SIZE-1) & MULT_13(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(8)(MULT_SIZE-1) & MULT_14(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(9)<=signed(MULT_13(9)(MULT_SIZE-1) & MULT_13(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(9)(MULT_SIZE-1) & MULT_14(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_8(0)<=signed(MULT_15(0)(MULT_SIZE-1) & MULT_15(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(0)(MULT_SIZE-1) & MULT_16(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(1)<=signed(MULT_15(1)(MULT_SIZE-1) & MULT_15(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(1)(MULT_SIZE-1) & MULT_16(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(2)<=signed(MULT_15(2)(MULT_SIZE-1) & MULT_15(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(2)(MULT_SIZE-1) & MULT_16(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(3)<=signed(MULT_15(3)(MULT_SIZE-1) & MULT_15(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(3)(MULT_SIZE-1) & MULT_16(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(4)<=signed(MULT_15(4)(MULT_SIZE-1) & MULT_15(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(4)(MULT_SIZE-1) & MULT_16(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(5)<=signed(MULT_15(5)(MULT_SIZE-1) & MULT_15(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(5)(MULT_SIZE-1) & MULT_16(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(6)<=signed(MULT_15(6)(MULT_SIZE-1) & MULT_15(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(6)(MULT_SIZE-1) & MULT_16(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(7)<=signed(MULT_15(7)(MULT_SIZE-1) & MULT_15(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(7)(MULT_SIZE-1) & MULT_16(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(8)<=signed(MULT_15(8)(MULT_SIZE-1) & MULT_15(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(8)(MULT_SIZE-1) & MULT_16(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(9)<=signed(MULT_15(9)(MULT_SIZE-1) & MULT_15(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(9)(MULT_SIZE-1) & MULT_16(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_9(0)<=signed(MULT_17(0)(MULT_SIZE-1) & MULT_17(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(0)(MULT_SIZE-1) & MULT_18(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(1)<=signed(MULT_17(1)(MULT_SIZE-1) & MULT_17(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(1)(MULT_SIZE-1) & MULT_18(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(2)<=signed(MULT_17(2)(MULT_SIZE-1) & MULT_17(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(2)(MULT_SIZE-1) & MULT_18(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(3)<=signed(MULT_17(3)(MULT_SIZE-1) & MULT_17(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(3)(MULT_SIZE-1) & MULT_18(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(4)<=signed(MULT_17(4)(MULT_SIZE-1) & MULT_17(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(4)(MULT_SIZE-1) & MULT_18(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(5)<=signed(MULT_17(5)(MULT_SIZE-1) & MULT_17(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(5)(MULT_SIZE-1) & MULT_18(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(6)<=signed(MULT_17(6)(MULT_SIZE-1) & MULT_17(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(6)(MULT_SIZE-1) & MULT_18(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(7)<=signed(MULT_17(7)(MULT_SIZE-1) & MULT_17(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(7)(MULT_SIZE-1) & MULT_18(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(8)<=signed(MULT_17(8)(MULT_SIZE-1) & MULT_17(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(8)(MULT_SIZE-1) & MULT_18(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(9)<=signed(MULT_17(9)(MULT_SIZE-1) & MULT_17(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(9)(MULT_SIZE-1) & MULT_18(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_10(0)<=signed(MULT_19(0)(MULT_SIZE-1) & MULT_19(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(0)(MULT_SIZE-1) & MULT_20(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(1)<=signed(MULT_19(1)(MULT_SIZE-1) & MULT_19(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(1)(MULT_SIZE-1) & MULT_20(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(2)<=signed(MULT_19(2)(MULT_SIZE-1) & MULT_19(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(2)(MULT_SIZE-1) & MULT_20(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(3)<=signed(MULT_19(3)(MULT_SIZE-1) & MULT_19(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(3)(MULT_SIZE-1) & MULT_20(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(4)<=signed(MULT_19(4)(MULT_SIZE-1) & MULT_19(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(4)(MULT_SIZE-1) & MULT_20(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(5)<=signed(MULT_19(5)(MULT_SIZE-1) & MULT_19(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(5)(MULT_SIZE-1) & MULT_20(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(6)<=signed(MULT_19(6)(MULT_SIZE-1) & MULT_19(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(6)(MULT_SIZE-1) & MULT_20(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(7)<=signed(MULT_19(7)(MULT_SIZE-1) & MULT_19(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(7)(MULT_SIZE-1) & MULT_20(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(8)<=signed(MULT_19(8)(MULT_SIZE-1) & MULT_19(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(8)(MULT_SIZE-1) & MULT_20(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(9)<=signed(MULT_19(9)(MULT_SIZE-1) & MULT_19(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(9)(MULT_SIZE-1) & MULT_20(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_11(0)<=signed(MULT_21(0)(MULT_SIZE-1) & MULT_21(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(0)(MULT_SIZE-1) & MULT_22(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(1)<=signed(MULT_21(1)(MULT_SIZE-1) & MULT_21(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(1)(MULT_SIZE-1) & MULT_22(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(2)<=signed(MULT_21(2)(MULT_SIZE-1) & MULT_21(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(2)(MULT_SIZE-1) & MULT_22(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(3)<=signed(MULT_21(3)(MULT_SIZE-1) & MULT_21(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(3)(MULT_SIZE-1) & MULT_22(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(4)<=signed(MULT_21(4)(MULT_SIZE-1) & MULT_21(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(4)(MULT_SIZE-1) & MULT_22(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(5)<=signed(MULT_21(5)(MULT_SIZE-1) & MULT_21(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(5)(MULT_SIZE-1) & MULT_22(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(6)<=signed(MULT_21(6)(MULT_SIZE-1) & MULT_21(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(6)(MULT_SIZE-1) & MULT_22(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(7)<=signed(MULT_21(7)(MULT_SIZE-1) & MULT_21(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(7)(MULT_SIZE-1) & MULT_22(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(8)<=signed(MULT_21(8)(MULT_SIZE-1) & MULT_21(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(8)(MULT_SIZE-1) & MULT_22(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(9)<=signed(MULT_21(9)(MULT_SIZE-1) & MULT_21(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(9)(MULT_SIZE-1) & MULT_22(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_12(0)<=signed(MULT_23(0)(MULT_SIZE-1) & MULT_23(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(0)(MULT_SIZE-1) & MULT_24(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(1)<=signed(MULT_23(1)(MULT_SIZE-1) & MULT_23(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(1)(MULT_SIZE-1) & MULT_24(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(2)<=signed(MULT_23(2)(MULT_SIZE-1) & MULT_23(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(2)(MULT_SIZE-1) & MULT_24(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(3)<=signed(MULT_23(3)(MULT_SIZE-1) & MULT_23(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(3)(MULT_SIZE-1) & MULT_24(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(4)<=signed(MULT_23(4)(MULT_SIZE-1) & MULT_23(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(4)(MULT_SIZE-1) & MULT_24(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(5)<=signed(MULT_23(5)(MULT_SIZE-1) & MULT_23(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(5)(MULT_SIZE-1) & MULT_24(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(6)<=signed(MULT_23(6)(MULT_SIZE-1) & MULT_23(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(6)(MULT_SIZE-1) & MULT_24(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(7)<=signed(MULT_23(7)(MULT_SIZE-1) & MULT_23(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(7)(MULT_SIZE-1) & MULT_24(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(8)<=signed(MULT_23(8)(MULT_SIZE-1) & MULT_23(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(8)(MULT_SIZE-1) & MULT_24(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(9)<=signed(MULT_23(9)(MULT_SIZE-1) & MULT_23(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(9)(MULT_SIZE-1) & MULT_24(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_13(0)<=signed(MULT_25(0)(MULT_SIZE-1) & MULT_25(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(0)(MULT_SIZE-1) & MULT_26(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(1)<=signed(MULT_25(1)(MULT_SIZE-1) & MULT_25(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(1)(MULT_SIZE-1) & MULT_26(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(2)<=signed(MULT_25(2)(MULT_SIZE-1) & MULT_25(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(2)(MULT_SIZE-1) & MULT_26(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(3)<=signed(MULT_25(3)(MULT_SIZE-1) & MULT_25(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(3)(MULT_SIZE-1) & MULT_26(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(4)<=signed(MULT_25(4)(MULT_SIZE-1) & MULT_25(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(4)(MULT_SIZE-1) & MULT_26(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(5)<=signed(MULT_25(5)(MULT_SIZE-1) & MULT_25(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(5)(MULT_SIZE-1) & MULT_26(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(6)<=signed(MULT_25(6)(MULT_SIZE-1) & MULT_25(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(6)(MULT_SIZE-1) & MULT_26(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(7)<=signed(MULT_25(7)(MULT_SIZE-1) & MULT_25(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(7)(MULT_SIZE-1) & MULT_26(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(8)<=signed(MULT_25(8)(MULT_SIZE-1) & MULT_25(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(8)(MULT_SIZE-1) & MULT_26(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(9)<=signed(MULT_25(9)(MULT_SIZE-1) & MULT_25(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(9)(MULT_SIZE-1) & MULT_26(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_14(0)<=signed(MULT_27(0)(MULT_SIZE-1) & MULT_27(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(0)(MULT_SIZE-1) & MULT_28(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(1)<=signed(MULT_27(1)(MULT_SIZE-1) & MULT_27(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(1)(MULT_SIZE-1) & MULT_28(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(2)<=signed(MULT_27(2)(MULT_SIZE-1) & MULT_27(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(2)(MULT_SIZE-1) & MULT_28(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(3)<=signed(MULT_27(3)(MULT_SIZE-1) & MULT_27(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(3)(MULT_SIZE-1) & MULT_28(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(4)<=signed(MULT_27(4)(MULT_SIZE-1) & MULT_27(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(4)(MULT_SIZE-1) & MULT_28(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(5)<=signed(MULT_27(5)(MULT_SIZE-1) & MULT_27(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(5)(MULT_SIZE-1) & MULT_28(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(6)<=signed(MULT_27(6)(MULT_SIZE-1) & MULT_27(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(6)(MULT_SIZE-1) & MULT_28(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(7)<=signed(MULT_27(7)(MULT_SIZE-1) & MULT_27(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(7)(MULT_SIZE-1) & MULT_28(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(8)<=signed(MULT_27(8)(MULT_SIZE-1) & MULT_27(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(8)(MULT_SIZE-1) & MULT_28(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(9)<=signed(MULT_27(9)(MULT_SIZE-1) & MULT_27(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(9)(MULT_SIZE-1) & MULT_28(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_15(0)<=signed(MULT_29(0)(MULT_SIZE-1) & MULT_29(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(0)(MULT_SIZE-1) & MULT_30(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(1)<=signed(MULT_29(1)(MULT_SIZE-1) & MULT_29(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(1)(MULT_SIZE-1) & MULT_30(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(2)<=signed(MULT_29(2)(MULT_SIZE-1) & MULT_29(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(2)(MULT_SIZE-1) & MULT_30(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(3)<=signed(MULT_29(3)(MULT_SIZE-1) & MULT_29(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(3)(MULT_SIZE-1) & MULT_30(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(4)<=signed(MULT_29(4)(MULT_SIZE-1) & MULT_29(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(4)(MULT_SIZE-1) & MULT_30(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(5)<=signed(MULT_29(5)(MULT_SIZE-1) & MULT_29(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(5)(MULT_SIZE-1) & MULT_30(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(6)<=signed(MULT_29(6)(MULT_SIZE-1) & MULT_29(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(6)(MULT_SIZE-1) & MULT_30(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(7)<=signed(MULT_29(7)(MULT_SIZE-1) & MULT_29(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(7)(MULT_SIZE-1) & MULT_30(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(8)<=signed(MULT_29(8)(MULT_SIZE-1) & MULT_29(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(8)(MULT_SIZE-1) & MULT_30(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(9)<=signed(MULT_29(9)(MULT_SIZE-1) & MULT_29(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(9)(MULT_SIZE-1) & MULT_30(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_16(0)<=signed(MULT_31(0)(MULT_SIZE-1) & MULT_31(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(0)(MULT_SIZE-1) & MULT_32(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(1)<=signed(MULT_31(1)(MULT_SIZE-1) & MULT_31(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(1)(MULT_SIZE-1) & MULT_32(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(2)<=signed(MULT_31(2)(MULT_SIZE-1) & MULT_31(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(2)(MULT_SIZE-1) & MULT_32(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(3)<=signed(MULT_31(3)(MULT_SIZE-1) & MULT_31(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(3)(MULT_SIZE-1) & MULT_32(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(4)<=signed(MULT_31(4)(MULT_SIZE-1) & MULT_31(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(4)(MULT_SIZE-1) & MULT_32(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(5)<=signed(MULT_31(5)(MULT_SIZE-1) & MULT_31(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(5)(MULT_SIZE-1) & MULT_32(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(6)<=signed(MULT_31(6)(MULT_SIZE-1) & MULT_31(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(6)(MULT_SIZE-1) & MULT_32(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(7)<=signed(MULT_31(7)(MULT_SIZE-1) & MULT_31(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(7)(MULT_SIZE-1) & MULT_32(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(8)<=signed(MULT_31(8)(MULT_SIZE-1) & MULT_31(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(8)(MULT_SIZE-1) & MULT_32(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(9)<=signed(MULT_31(9)(MULT_SIZE-1) & MULT_31(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(9)(MULT_SIZE-1) & MULT_32(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_17(0)<=signed(MULT_33(0)(MULT_SIZE-1) & MULT_33(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(0)(MULT_SIZE-1) & MULT_34(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(1)<=signed(MULT_33(1)(MULT_SIZE-1) & MULT_33(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(1)(MULT_SIZE-1) & MULT_34(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(2)<=signed(MULT_33(2)(MULT_SIZE-1) & MULT_33(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(2)(MULT_SIZE-1) & MULT_34(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(3)<=signed(MULT_33(3)(MULT_SIZE-1) & MULT_33(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(3)(MULT_SIZE-1) & MULT_34(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(4)<=signed(MULT_33(4)(MULT_SIZE-1) & MULT_33(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(4)(MULT_SIZE-1) & MULT_34(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(5)<=signed(MULT_33(5)(MULT_SIZE-1) & MULT_33(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(5)(MULT_SIZE-1) & MULT_34(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(6)<=signed(MULT_33(6)(MULT_SIZE-1) & MULT_33(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(6)(MULT_SIZE-1) & MULT_34(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(7)<=signed(MULT_33(7)(MULT_SIZE-1) & MULT_33(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(7)(MULT_SIZE-1) & MULT_34(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(8)<=signed(MULT_33(8)(MULT_SIZE-1) & MULT_33(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(8)(MULT_SIZE-1) & MULT_34(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(9)<=signed(MULT_33(9)(MULT_SIZE-1) & MULT_33(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(9)(MULT_SIZE-1) & MULT_34(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_18(0)<=signed(MULT_35(0)(MULT_SIZE-1) & MULT_35(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(0)(MULT_SIZE-1) & MULT_36(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(1)<=signed(MULT_35(1)(MULT_SIZE-1) & MULT_35(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(1)(MULT_SIZE-1) & MULT_36(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(2)<=signed(MULT_35(2)(MULT_SIZE-1) & MULT_35(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(2)(MULT_SIZE-1) & MULT_36(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(3)<=signed(MULT_35(3)(MULT_SIZE-1) & MULT_35(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(3)(MULT_SIZE-1) & MULT_36(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(4)<=signed(MULT_35(4)(MULT_SIZE-1) & MULT_35(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(4)(MULT_SIZE-1) & MULT_36(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(5)<=signed(MULT_35(5)(MULT_SIZE-1) & MULT_35(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(5)(MULT_SIZE-1) & MULT_36(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(6)<=signed(MULT_35(6)(MULT_SIZE-1) & MULT_35(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(6)(MULT_SIZE-1) & MULT_36(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(7)<=signed(MULT_35(7)(MULT_SIZE-1) & MULT_35(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(7)(MULT_SIZE-1) & MULT_36(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(8)<=signed(MULT_35(8)(MULT_SIZE-1) & MULT_35(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(8)(MULT_SIZE-1) & MULT_36(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(9)<=signed(MULT_35(9)(MULT_SIZE-1) & MULT_35(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(9)(MULT_SIZE-1) & MULT_36(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_19(0)<=signed(MULT_37(0)(MULT_SIZE-1) & MULT_37(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(0)(MULT_SIZE-1) & MULT_38(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(1)<=signed(MULT_37(1)(MULT_SIZE-1) & MULT_37(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(1)(MULT_SIZE-1) & MULT_38(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(2)<=signed(MULT_37(2)(MULT_SIZE-1) & MULT_37(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(2)(MULT_SIZE-1) & MULT_38(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(3)<=signed(MULT_37(3)(MULT_SIZE-1) & MULT_37(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(3)(MULT_SIZE-1) & MULT_38(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(4)<=signed(MULT_37(4)(MULT_SIZE-1) & MULT_37(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(4)(MULT_SIZE-1) & MULT_38(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(5)<=signed(MULT_37(5)(MULT_SIZE-1) & MULT_37(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(5)(MULT_SIZE-1) & MULT_38(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(6)<=signed(MULT_37(6)(MULT_SIZE-1) & MULT_37(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(6)(MULT_SIZE-1) & MULT_38(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(7)<=signed(MULT_37(7)(MULT_SIZE-1) & MULT_37(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(7)(MULT_SIZE-1) & MULT_38(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(8)<=signed(MULT_37(8)(MULT_SIZE-1) & MULT_37(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(8)(MULT_SIZE-1) & MULT_38(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(9)<=signed(MULT_37(9)(MULT_SIZE-1) & MULT_37(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(9)(MULT_SIZE-1) & MULT_38(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_20(0)<=signed(MULT_39(0)(MULT_SIZE-1) & MULT_39(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(0)(MULT_SIZE-1) & MULT_40(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(1)<=signed(MULT_39(1)(MULT_SIZE-1) & MULT_39(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(1)(MULT_SIZE-1) & MULT_40(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(2)<=signed(MULT_39(2)(MULT_SIZE-1) & MULT_39(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(2)(MULT_SIZE-1) & MULT_40(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(3)<=signed(MULT_39(3)(MULT_SIZE-1) & MULT_39(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(3)(MULT_SIZE-1) & MULT_40(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(4)<=signed(MULT_39(4)(MULT_SIZE-1) & MULT_39(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(4)(MULT_SIZE-1) & MULT_40(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(5)<=signed(MULT_39(5)(MULT_SIZE-1) & MULT_39(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(5)(MULT_SIZE-1) & MULT_40(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(6)<=signed(MULT_39(6)(MULT_SIZE-1) & MULT_39(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(6)(MULT_SIZE-1) & MULT_40(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(7)<=signed(MULT_39(7)(MULT_SIZE-1) & MULT_39(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(7)(MULT_SIZE-1) & MULT_40(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(8)<=signed(MULT_39(8)(MULT_SIZE-1) & MULT_39(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(8)(MULT_SIZE-1) & MULT_40(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(9)<=signed(MULT_39(9)(MULT_SIZE-1) & MULT_39(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(9)(MULT_SIZE-1) & MULT_40(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_21(0)<=signed(MULT_41(0)(MULT_SIZE-1) & MULT_41(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(0)(MULT_SIZE-1) & MULT_42(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(1)<=signed(MULT_41(1)(MULT_SIZE-1) & MULT_41(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(1)(MULT_SIZE-1) & MULT_42(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(2)<=signed(MULT_41(2)(MULT_SIZE-1) & MULT_41(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(2)(MULT_SIZE-1) & MULT_42(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(3)<=signed(MULT_41(3)(MULT_SIZE-1) & MULT_41(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(3)(MULT_SIZE-1) & MULT_42(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(4)<=signed(MULT_41(4)(MULT_SIZE-1) & MULT_41(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(4)(MULT_SIZE-1) & MULT_42(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(5)<=signed(MULT_41(5)(MULT_SIZE-1) & MULT_41(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(5)(MULT_SIZE-1) & MULT_42(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(6)<=signed(MULT_41(6)(MULT_SIZE-1) & MULT_41(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(6)(MULT_SIZE-1) & MULT_42(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(7)<=signed(MULT_41(7)(MULT_SIZE-1) & MULT_41(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(7)(MULT_SIZE-1) & MULT_42(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(8)<=signed(MULT_41(8)(MULT_SIZE-1) & MULT_41(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(8)(MULT_SIZE-1) & MULT_42(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(9)<=signed(MULT_41(9)(MULT_SIZE-1) & MULT_41(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(9)(MULT_SIZE-1) & MULT_42(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_22(0)<=signed(MULT_43(0)(MULT_SIZE-1) & MULT_43(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(0)(MULT_SIZE-1) & MULT_44(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(1)<=signed(MULT_43(1)(MULT_SIZE-1) & MULT_43(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(1)(MULT_SIZE-1) & MULT_44(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(2)<=signed(MULT_43(2)(MULT_SIZE-1) & MULT_43(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(2)(MULT_SIZE-1) & MULT_44(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(3)<=signed(MULT_43(3)(MULT_SIZE-1) & MULT_43(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(3)(MULT_SIZE-1) & MULT_44(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(4)<=signed(MULT_43(4)(MULT_SIZE-1) & MULT_43(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(4)(MULT_SIZE-1) & MULT_44(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(5)<=signed(MULT_43(5)(MULT_SIZE-1) & MULT_43(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(5)(MULT_SIZE-1) & MULT_44(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(6)<=signed(MULT_43(6)(MULT_SIZE-1) & MULT_43(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(6)(MULT_SIZE-1) & MULT_44(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(7)<=signed(MULT_43(7)(MULT_SIZE-1) & MULT_43(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(7)(MULT_SIZE-1) & MULT_44(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(8)<=signed(MULT_43(8)(MULT_SIZE-1) & MULT_43(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(8)(MULT_SIZE-1) & MULT_44(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(9)<=signed(MULT_43(9)(MULT_SIZE-1) & MULT_43(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(9)(MULT_SIZE-1) & MULT_44(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_23(0)<=signed(MULT_45(0)(MULT_SIZE-1) & MULT_45(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(0)(MULT_SIZE-1) & MULT_46(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(1)<=signed(MULT_45(1)(MULT_SIZE-1) & MULT_45(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(1)(MULT_SIZE-1) & MULT_46(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(2)<=signed(MULT_45(2)(MULT_SIZE-1) & MULT_45(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(2)(MULT_SIZE-1) & MULT_46(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(3)<=signed(MULT_45(3)(MULT_SIZE-1) & MULT_45(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(3)(MULT_SIZE-1) & MULT_46(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(4)<=signed(MULT_45(4)(MULT_SIZE-1) & MULT_45(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(4)(MULT_SIZE-1) & MULT_46(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(5)<=signed(MULT_45(5)(MULT_SIZE-1) & MULT_45(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(5)(MULT_SIZE-1) & MULT_46(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(6)<=signed(MULT_45(6)(MULT_SIZE-1) & MULT_45(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(6)(MULT_SIZE-1) & MULT_46(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(7)<=signed(MULT_45(7)(MULT_SIZE-1) & MULT_45(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(7)(MULT_SIZE-1) & MULT_46(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(8)<=signed(MULT_45(8)(MULT_SIZE-1) & MULT_45(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(8)(MULT_SIZE-1) & MULT_46(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(9)<=signed(MULT_45(9)(MULT_SIZE-1) & MULT_45(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(9)(MULT_SIZE-1) & MULT_46(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_24(0)<=signed(MULT_47(0)(MULT_SIZE-1) & MULT_47(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(0)(MULT_SIZE-1) & MULT_48(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(1)<=signed(MULT_47(1)(MULT_SIZE-1) & MULT_47(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(1)(MULT_SIZE-1) & MULT_48(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(2)<=signed(MULT_47(2)(MULT_SIZE-1) & MULT_47(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(2)(MULT_SIZE-1) & MULT_48(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(3)<=signed(MULT_47(3)(MULT_SIZE-1) & MULT_47(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(3)(MULT_SIZE-1) & MULT_48(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(4)<=signed(MULT_47(4)(MULT_SIZE-1) & MULT_47(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(4)(MULT_SIZE-1) & MULT_48(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(5)<=signed(MULT_47(5)(MULT_SIZE-1) & MULT_47(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(5)(MULT_SIZE-1) & MULT_48(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(6)<=signed(MULT_47(6)(MULT_SIZE-1) & MULT_47(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(6)(MULT_SIZE-1) & MULT_48(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(7)<=signed(MULT_47(7)(MULT_SIZE-1) & MULT_47(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(7)(MULT_SIZE-1) & MULT_48(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(8)<=signed(MULT_47(8)(MULT_SIZE-1) & MULT_47(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(8)(MULT_SIZE-1) & MULT_48(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(9)<=signed(MULT_47(9)(MULT_SIZE-1) & MULT_47(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(9)(MULT_SIZE-1) & MULT_48(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_25(0)<=signed(MULT_49(0)(MULT_SIZE-1) & MULT_49(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(0)(MULT_SIZE-1) & MULT_50(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(1)<=signed(MULT_49(1)(MULT_SIZE-1) & MULT_49(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(1)(MULT_SIZE-1) & MULT_50(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(2)<=signed(MULT_49(2)(MULT_SIZE-1) & MULT_49(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(2)(MULT_SIZE-1) & MULT_50(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(3)<=signed(MULT_49(3)(MULT_SIZE-1) & MULT_49(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(3)(MULT_SIZE-1) & MULT_50(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(4)<=signed(MULT_49(4)(MULT_SIZE-1) & MULT_49(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(4)(MULT_SIZE-1) & MULT_50(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(5)<=signed(MULT_49(5)(MULT_SIZE-1) & MULT_49(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(5)(MULT_SIZE-1) & MULT_50(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(6)<=signed(MULT_49(6)(MULT_SIZE-1) & MULT_49(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(6)(MULT_SIZE-1) & MULT_50(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(7)<=signed(MULT_49(7)(MULT_SIZE-1) & MULT_49(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(7)(MULT_SIZE-1) & MULT_50(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(8)<=signed(MULT_49(8)(MULT_SIZE-1) & MULT_49(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(8)(MULT_SIZE-1) & MULT_50(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(9)<=signed(MULT_49(9)(MULT_SIZE-1) & MULT_49(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(9)(MULT_SIZE-1) & MULT_50(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_26(0)<=signed(MULT_51(0)(MULT_SIZE-1) & MULT_51(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(0)(MULT_SIZE-1) & MULT_52(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(1)<=signed(MULT_51(1)(MULT_SIZE-1) & MULT_51(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(1)(MULT_SIZE-1) & MULT_52(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(2)<=signed(MULT_51(2)(MULT_SIZE-1) & MULT_51(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(2)(MULT_SIZE-1) & MULT_52(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(3)<=signed(MULT_51(3)(MULT_SIZE-1) & MULT_51(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(3)(MULT_SIZE-1) & MULT_52(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(4)<=signed(MULT_51(4)(MULT_SIZE-1) & MULT_51(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(4)(MULT_SIZE-1) & MULT_52(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(5)<=signed(MULT_51(5)(MULT_SIZE-1) & MULT_51(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(5)(MULT_SIZE-1) & MULT_52(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(6)<=signed(MULT_51(6)(MULT_SIZE-1) & MULT_51(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(6)(MULT_SIZE-1) & MULT_52(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(7)<=signed(MULT_51(7)(MULT_SIZE-1) & MULT_51(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(7)(MULT_SIZE-1) & MULT_52(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(8)<=signed(MULT_51(8)(MULT_SIZE-1) & MULT_51(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(8)(MULT_SIZE-1) & MULT_52(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(9)<=signed(MULT_51(9)(MULT_SIZE-1) & MULT_51(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(9)(MULT_SIZE-1) & MULT_52(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_27(0)<=signed(MULT_53(0)(MULT_SIZE-1) & MULT_53(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(0)(MULT_SIZE-1) & MULT_54(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(1)<=signed(MULT_53(1)(MULT_SIZE-1) & MULT_53(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(1)(MULT_SIZE-1) & MULT_54(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(2)<=signed(MULT_53(2)(MULT_SIZE-1) & MULT_53(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(2)(MULT_SIZE-1) & MULT_54(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(3)<=signed(MULT_53(3)(MULT_SIZE-1) & MULT_53(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(3)(MULT_SIZE-1) & MULT_54(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(4)<=signed(MULT_53(4)(MULT_SIZE-1) & MULT_53(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(4)(MULT_SIZE-1) & MULT_54(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(5)<=signed(MULT_53(5)(MULT_SIZE-1) & MULT_53(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(5)(MULT_SIZE-1) & MULT_54(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(6)<=signed(MULT_53(6)(MULT_SIZE-1) & MULT_53(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(6)(MULT_SIZE-1) & MULT_54(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(7)<=signed(MULT_53(7)(MULT_SIZE-1) & MULT_53(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(7)(MULT_SIZE-1) & MULT_54(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(8)<=signed(MULT_53(8)(MULT_SIZE-1) & MULT_53(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(8)(MULT_SIZE-1) & MULT_54(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(9)<=signed(MULT_53(9)(MULT_SIZE-1) & MULT_53(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(9)(MULT_SIZE-1) & MULT_54(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_28(0)<=signed(MULT_55(0)(MULT_SIZE-1) & MULT_55(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(0)(MULT_SIZE-1) & MULT_56(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(1)<=signed(MULT_55(1)(MULT_SIZE-1) & MULT_55(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(1)(MULT_SIZE-1) & MULT_56(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(2)<=signed(MULT_55(2)(MULT_SIZE-1) & MULT_55(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(2)(MULT_SIZE-1) & MULT_56(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(3)<=signed(MULT_55(3)(MULT_SIZE-1) & MULT_55(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(3)(MULT_SIZE-1) & MULT_56(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(4)<=signed(MULT_55(4)(MULT_SIZE-1) & MULT_55(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(4)(MULT_SIZE-1) & MULT_56(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(5)<=signed(MULT_55(5)(MULT_SIZE-1) & MULT_55(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(5)(MULT_SIZE-1) & MULT_56(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(6)<=signed(MULT_55(6)(MULT_SIZE-1) & MULT_55(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(6)(MULT_SIZE-1) & MULT_56(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(7)<=signed(MULT_55(7)(MULT_SIZE-1) & MULT_55(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(7)(MULT_SIZE-1) & MULT_56(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(8)<=signed(MULT_55(8)(MULT_SIZE-1) & MULT_55(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(8)(MULT_SIZE-1) & MULT_56(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(9)<=signed(MULT_55(9)(MULT_SIZE-1) & MULT_55(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(9)(MULT_SIZE-1) & MULT_56(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_29(0)<=signed(MULT_57(0)(MULT_SIZE-1) & MULT_57(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(0)(MULT_SIZE-1) & MULT_58(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(1)<=signed(MULT_57(1)(MULT_SIZE-1) & MULT_57(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(1)(MULT_SIZE-1) & MULT_58(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(2)<=signed(MULT_57(2)(MULT_SIZE-1) & MULT_57(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(2)(MULT_SIZE-1) & MULT_58(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(3)<=signed(MULT_57(3)(MULT_SIZE-1) & MULT_57(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(3)(MULT_SIZE-1) & MULT_58(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(4)<=signed(MULT_57(4)(MULT_SIZE-1) & MULT_57(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(4)(MULT_SIZE-1) & MULT_58(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(5)<=signed(MULT_57(5)(MULT_SIZE-1) & MULT_57(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(5)(MULT_SIZE-1) & MULT_58(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(6)<=signed(MULT_57(6)(MULT_SIZE-1) & MULT_57(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(6)(MULT_SIZE-1) & MULT_58(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(7)<=signed(MULT_57(7)(MULT_SIZE-1) & MULT_57(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(7)(MULT_SIZE-1) & MULT_58(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(8)<=signed(MULT_57(8)(MULT_SIZE-1) & MULT_57(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(8)(MULT_SIZE-1) & MULT_58(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(9)<=signed(MULT_57(9)(MULT_SIZE-1) & MULT_57(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(9)(MULT_SIZE-1) & MULT_58(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_30(0)<=signed(MULT_59(0)(MULT_SIZE-1) & MULT_59(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(0)(MULT_SIZE-1) & MULT_60(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(1)<=signed(MULT_59(1)(MULT_SIZE-1) & MULT_59(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(1)(MULT_SIZE-1) & MULT_60(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(2)<=signed(MULT_59(2)(MULT_SIZE-1) & MULT_59(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(2)(MULT_SIZE-1) & MULT_60(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(3)<=signed(MULT_59(3)(MULT_SIZE-1) & MULT_59(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(3)(MULT_SIZE-1) & MULT_60(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(4)<=signed(MULT_59(4)(MULT_SIZE-1) & MULT_59(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(4)(MULT_SIZE-1) & MULT_60(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(5)<=signed(MULT_59(5)(MULT_SIZE-1) & MULT_59(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(5)(MULT_SIZE-1) & MULT_60(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(6)<=signed(MULT_59(6)(MULT_SIZE-1) & MULT_59(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(6)(MULT_SIZE-1) & MULT_60(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(7)<=signed(MULT_59(7)(MULT_SIZE-1) & MULT_59(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(7)(MULT_SIZE-1) & MULT_60(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(8)<=signed(MULT_59(8)(MULT_SIZE-1) & MULT_59(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(8)(MULT_SIZE-1) & MULT_60(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(9)<=signed(MULT_59(9)(MULT_SIZE-1) & MULT_59(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(9)(MULT_SIZE-1) & MULT_60(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_31(0)<=signed(MULT_61(0)(MULT_SIZE-1) & MULT_61(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(0)(MULT_SIZE-1) & MULT_62(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(1)<=signed(MULT_61(1)(MULT_SIZE-1) & MULT_61(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(1)(MULT_SIZE-1) & MULT_62(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(2)<=signed(MULT_61(2)(MULT_SIZE-1) & MULT_61(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(2)(MULT_SIZE-1) & MULT_62(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(3)<=signed(MULT_61(3)(MULT_SIZE-1) & MULT_61(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(3)(MULT_SIZE-1) & MULT_62(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(4)<=signed(MULT_61(4)(MULT_SIZE-1) & MULT_61(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(4)(MULT_SIZE-1) & MULT_62(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(5)<=signed(MULT_61(5)(MULT_SIZE-1) & MULT_61(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(5)(MULT_SIZE-1) & MULT_62(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(6)<=signed(MULT_61(6)(MULT_SIZE-1) & MULT_61(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(6)(MULT_SIZE-1) & MULT_62(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(7)<=signed(MULT_61(7)(MULT_SIZE-1) & MULT_61(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(7)(MULT_SIZE-1) & MULT_62(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(8)<=signed(MULT_61(8)(MULT_SIZE-1) & MULT_61(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(8)(MULT_SIZE-1) & MULT_62(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(9)<=signed(MULT_61(9)(MULT_SIZE-1) & MULT_61(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(9)(MULT_SIZE-1) & MULT_62(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_32(0)<=signed(MULT_63(0)(MULT_SIZE-1) & MULT_63(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(0)(MULT_SIZE-1) & MULT_64(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(1)<=signed(MULT_63(1)(MULT_SIZE-1) & MULT_63(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(1)(MULT_SIZE-1) & MULT_64(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(2)<=signed(MULT_63(2)(MULT_SIZE-1) & MULT_63(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(2)(MULT_SIZE-1) & MULT_64(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(3)<=signed(MULT_63(3)(MULT_SIZE-1) & MULT_63(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(3)(MULT_SIZE-1) & MULT_64(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(4)<=signed(MULT_63(4)(MULT_SIZE-1) & MULT_63(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(4)(MULT_SIZE-1) & MULT_64(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(5)<=signed(MULT_63(5)(MULT_SIZE-1) & MULT_63(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(5)(MULT_SIZE-1) & MULT_64(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(6)<=signed(MULT_63(6)(MULT_SIZE-1) & MULT_63(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(6)(MULT_SIZE-1) & MULT_64(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(7)<=signed(MULT_63(7)(MULT_SIZE-1) & MULT_63(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(7)(MULT_SIZE-1) & MULT_64(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(8)<=signed(MULT_63(8)(MULT_SIZE-1) & MULT_63(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(8)(MULT_SIZE-1) & MULT_64(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(9)<=signed(MULT_63(9)(MULT_SIZE-1) & MULT_63(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(9)(MULT_SIZE-1) & MULT_64(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_33(0)<=signed(MULT_65(0)(MULT_SIZE-1) & MULT_65(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(0)(MULT_SIZE-1) & MULT_66(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(1)<=signed(MULT_65(1)(MULT_SIZE-1) & MULT_65(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(1)(MULT_SIZE-1) & MULT_66(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(2)<=signed(MULT_65(2)(MULT_SIZE-1) & MULT_65(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(2)(MULT_SIZE-1) & MULT_66(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(3)<=signed(MULT_65(3)(MULT_SIZE-1) & MULT_65(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(3)(MULT_SIZE-1) & MULT_66(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(4)<=signed(MULT_65(4)(MULT_SIZE-1) & MULT_65(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(4)(MULT_SIZE-1) & MULT_66(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(5)<=signed(MULT_65(5)(MULT_SIZE-1) & MULT_65(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(5)(MULT_SIZE-1) & MULT_66(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(6)<=signed(MULT_65(6)(MULT_SIZE-1) & MULT_65(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(6)(MULT_SIZE-1) & MULT_66(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(7)<=signed(MULT_65(7)(MULT_SIZE-1) & MULT_65(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(7)(MULT_SIZE-1) & MULT_66(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(8)<=signed(MULT_65(8)(MULT_SIZE-1) & MULT_65(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(8)(MULT_SIZE-1) & MULT_66(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(9)<=signed(MULT_65(9)(MULT_SIZE-1) & MULT_65(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(9)(MULT_SIZE-1) & MULT_66(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_34(0)<=signed(MULT_67(0)(MULT_SIZE-1) & MULT_67(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(0)(MULT_SIZE-1) & MULT_68(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(1)<=signed(MULT_67(1)(MULT_SIZE-1) & MULT_67(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(1)(MULT_SIZE-1) & MULT_68(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(2)<=signed(MULT_67(2)(MULT_SIZE-1) & MULT_67(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(2)(MULT_SIZE-1) & MULT_68(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(3)<=signed(MULT_67(3)(MULT_SIZE-1) & MULT_67(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(3)(MULT_SIZE-1) & MULT_68(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(4)<=signed(MULT_67(4)(MULT_SIZE-1) & MULT_67(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(4)(MULT_SIZE-1) & MULT_68(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(5)<=signed(MULT_67(5)(MULT_SIZE-1) & MULT_67(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(5)(MULT_SIZE-1) & MULT_68(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(6)<=signed(MULT_67(6)(MULT_SIZE-1) & MULT_67(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(6)(MULT_SIZE-1) & MULT_68(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(7)<=signed(MULT_67(7)(MULT_SIZE-1) & MULT_67(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(7)(MULT_SIZE-1) & MULT_68(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(8)<=signed(MULT_67(8)(MULT_SIZE-1) & MULT_67(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(8)(MULT_SIZE-1) & MULT_68(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(9)<=signed(MULT_67(9)(MULT_SIZE-1) & MULT_67(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(9)(MULT_SIZE-1) & MULT_68(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_35(0)<=signed(MULT_69(0)(MULT_SIZE-1) & MULT_69(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(0)(MULT_SIZE-1) & MULT_70(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(1)<=signed(MULT_69(1)(MULT_SIZE-1) & MULT_69(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(1)(MULT_SIZE-1) & MULT_70(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(2)<=signed(MULT_69(2)(MULT_SIZE-1) & MULT_69(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(2)(MULT_SIZE-1) & MULT_70(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(3)<=signed(MULT_69(3)(MULT_SIZE-1) & MULT_69(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(3)(MULT_SIZE-1) & MULT_70(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(4)<=signed(MULT_69(4)(MULT_SIZE-1) & MULT_69(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(4)(MULT_SIZE-1) & MULT_70(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(5)<=signed(MULT_69(5)(MULT_SIZE-1) & MULT_69(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(5)(MULT_SIZE-1) & MULT_70(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(6)<=signed(MULT_69(6)(MULT_SIZE-1) & MULT_69(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(6)(MULT_SIZE-1) & MULT_70(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(7)<=signed(MULT_69(7)(MULT_SIZE-1) & MULT_69(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(7)(MULT_SIZE-1) & MULT_70(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(8)<=signed(MULT_69(8)(MULT_SIZE-1) & MULT_69(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(8)(MULT_SIZE-1) & MULT_70(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(9)<=signed(MULT_69(9)(MULT_SIZE-1) & MULT_69(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(9)(MULT_SIZE-1) & MULT_70(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_36(0)<=signed(MULT_71(0)(MULT_SIZE-1) & MULT_71(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(0)(MULT_SIZE-1) & MULT_72(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(1)<=signed(MULT_71(1)(MULT_SIZE-1) & MULT_71(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(1)(MULT_SIZE-1) & MULT_72(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(2)<=signed(MULT_71(2)(MULT_SIZE-1) & MULT_71(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(2)(MULT_SIZE-1) & MULT_72(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(3)<=signed(MULT_71(3)(MULT_SIZE-1) & MULT_71(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(3)(MULT_SIZE-1) & MULT_72(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(4)<=signed(MULT_71(4)(MULT_SIZE-1) & MULT_71(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(4)(MULT_SIZE-1) & MULT_72(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(5)<=signed(MULT_71(5)(MULT_SIZE-1) & MULT_71(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(5)(MULT_SIZE-1) & MULT_72(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(6)<=signed(MULT_71(6)(MULT_SIZE-1) & MULT_71(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(6)(MULT_SIZE-1) & MULT_72(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(7)<=signed(MULT_71(7)(MULT_SIZE-1) & MULT_71(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(7)(MULT_SIZE-1) & MULT_72(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(8)<=signed(MULT_71(8)(MULT_SIZE-1) & MULT_71(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(8)(MULT_SIZE-1) & MULT_72(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(9)<=signed(MULT_71(9)(MULT_SIZE-1) & MULT_71(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(9)(MULT_SIZE-1) & MULT_72(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_37(0)<=signed(MULT_73(0)(MULT_SIZE-1) & MULT_73(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(0)(MULT_SIZE-1) & MULT_74(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(1)<=signed(MULT_73(1)(MULT_SIZE-1) & MULT_73(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(1)(MULT_SIZE-1) & MULT_74(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(2)<=signed(MULT_73(2)(MULT_SIZE-1) & MULT_73(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(2)(MULT_SIZE-1) & MULT_74(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(3)<=signed(MULT_73(3)(MULT_SIZE-1) & MULT_73(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(3)(MULT_SIZE-1) & MULT_74(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(4)<=signed(MULT_73(4)(MULT_SIZE-1) & MULT_73(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(4)(MULT_SIZE-1) & MULT_74(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(5)<=signed(MULT_73(5)(MULT_SIZE-1) & MULT_73(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(5)(MULT_SIZE-1) & MULT_74(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(6)<=signed(MULT_73(6)(MULT_SIZE-1) & MULT_73(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(6)(MULT_SIZE-1) & MULT_74(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(7)<=signed(MULT_73(7)(MULT_SIZE-1) & MULT_73(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(7)(MULT_SIZE-1) & MULT_74(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(8)<=signed(MULT_73(8)(MULT_SIZE-1) & MULT_73(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(8)(MULT_SIZE-1) & MULT_74(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(9)<=signed(MULT_73(9)(MULT_SIZE-1) & MULT_73(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(9)(MULT_SIZE-1) & MULT_74(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_38(0)<=signed(MULT_75(0)(MULT_SIZE-1) & MULT_75(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(0)(MULT_SIZE-1) & MULT_76(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(1)<=signed(MULT_75(1)(MULT_SIZE-1) & MULT_75(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(1)(MULT_SIZE-1) & MULT_76(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(2)<=signed(MULT_75(2)(MULT_SIZE-1) & MULT_75(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(2)(MULT_SIZE-1) & MULT_76(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(3)<=signed(MULT_75(3)(MULT_SIZE-1) & MULT_75(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(3)(MULT_SIZE-1) & MULT_76(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(4)<=signed(MULT_75(4)(MULT_SIZE-1) & MULT_75(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(4)(MULT_SIZE-1) & MULT_76(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(5)<=signed(MULT_75(5)(MULT_SIZE-1) & MULT_75(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(5)(MULT_SIZE-1) & MULT_76(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(6)<=signed(MULT_75(6)(MULT_SIZE-1) & MULT_75(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(6)(MULT_SIZE-1) & MULT_76(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(7)<=signed(MULT_75(7)(MULT_SIZE-1) & MULT_75(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(7)(MULT_SIZE-1) & MULT_76(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(8)<=signed(MULT_75(8)(MULT_SIZE-1) & MULT_75(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(8)(MULT_SIZE-1) & MULT_76(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(9)<=signed(MULT_75(9)(MULT_SIZE-1) & MULT_75(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(9)(MULT_SIZE-1) & MULT_76(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_39(0)<=signed(MULT_77(0)(MULT_SIZE-1) & MULT_77(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(0)(MULT_SIZE-1) & MULT_78(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(1)<=signed(MULT_77(1)(MULT_SIZE-1) & MULT_77(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(1)(MULT_SIZE-1) & MULT_78(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(2)<=signed(MULT_77(2)(MULT_SIZE-1) & MULT_77(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(2)(MULT_SIZE-1) & MULT_78(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(3)<=signed(MULT_77(3)(MULT_SIZE-1) & MULT_77(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(3)(MULT_SIZE-1) & MULT_78(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(4)<=signed(MULT_77(4)(MULT_SIZE-1) & MULT_77(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(4)(MULT_SIZE-1) & MULT_78(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(5)<=signed(MULT_77(5)(MULT_SIZE-1) & MULT_77(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(5)(MULT_SIZE-1) & MULT_78(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(6)<=signed(MULT_77(6)(MULT_SIZE-1) & MULT_77(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(6)(MULT_SIZE-1) & MULT_78(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(7)<=signed(MULT_77(7)(MULT_SIZE-1) & MULT_77(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(7)(MULT_SIZE-1) & MULT_78(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(8)<=signed(MULT_77(8)(MULT_SIZE-1) & MULT_77(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(8)(MULT_SIZE-1) & MULT_78(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(9)<=signed(MULT_77(9)(MULT_SIZE-1) & MULT_77(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(9)(MULT_SIZE-1) & MULT_78(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_40(0)<=signed(MULT_79(0)(MULT_SIZE-1) & MULT_79(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(0)(MULT_SIZE-1) & MULT_80(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(1)<=signed(MULT_79(1)(MULT_SIZE-1) & MULT_79(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(1)(MULT_SIZE-1) & MULT_80(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(2)<=signed(MULT_79(2)(MULT_SIZE-1) & MULT_79(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(2)(MULT_SIZE-1) & MULT_80(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(3)<=signed(MULT_79(3)(MULT_SIZE-1) & MULT_79(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(3)(MULT_SIZE-1) & MULT_80(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(4)<=signed(MULT_79(4)(MULT_SIZE-1) & MULT_79(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(4)(MULT_SIZE-1) & MULT_80(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(5)<=signed(MULT_79(5)(MULT_SIZE-1) & MULT_79(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(5)(MULT_SIZE-1) & MULT_80(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(6)<=signed(MULT_79(6)(MULT_SIZE-1) & MULT_79(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(6)(MULT_SIZE-1) & MULT_80(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(7)<=signed(MULT_79(7)(MULT_SIZE-1) & MULT_79(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(7)(MULT_SIZE-1) & MULT_80(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(8)<=signed(MULT_79(8)(MULT_SIZE-1) & MULT_79(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(8)(MULT_SIZE-1) & MULT_80(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(9)<=signed(MULT_79(9)(MULT_SIZE-1) & MULT_79(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(9)(MULT_SIZE-1) & MULT_80(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_41(0)<=signed(MULT_81(0)(MULT_SIZE-1) & MULT_81(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(0)(MULT_SIZE-1) & MULT_82(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(1)<=signed(MULT_81(1)(MULT_SIZE-1) & MULT_81(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(1)(MULT_SIZE-1) & MULT_82(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(2)<=signed(MULT_81(2)(MULT_SIZE-1) & MULT_81(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(2)(MULT_SIZE-1) & MULT_82(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(3)<=signed(MULT_81(3)(MULT_SIZE-1) & MULT_81(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(3)(MULT_SIZE-1) & MULT_82(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(4)<=signed(MULT_81(4)(MULT_SIZE-1) & MULT_81(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(4)(MULT_SIZE-1) & MULT_82(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(5)<=signed(MULT_81(5)(MULT_SIZE-1) & MULT_81(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(5)(MULT_SIZE-1) & MULT_82(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(6)<=signed(MULT_81(6)(MULT_SIZE-1) & MULT_81(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(6)(MULT_SIZE-1) & MULT_82(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(7)<=signed(MULT_81(7)(MULT_SIZE-1) & MULT_81(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(7)(MULT_SIZE-1) & MULT_82(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(8)<=signed(MULT_81(8)(MULT_SIZE-1) & MULT_81(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(8)(MULT_SIZE-1) & MULT_82(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(9)<=signed(MULT_81(9)(MULT_SIZE-1) & MULT_81(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(9)(MULT_SIZE-1) & MULT_82(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_42(0)<=signed(MULT_83(0)(MULT_SIZE-1) & MULT_83(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(0)(MULT_SIZE-1) & MULT_84(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(1)<=signed(MULT_83(1)(MULT_SIZE-1) & MULT_83(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(1)(MULT_SIZE-1) & MULT_84(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(2)<=signed(MULT_83(2)(MULT_SIZE-1) & MULT_83(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(2)(MULT_SIZE-1) & MULT_84(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(3)<=signed(MULT_83(3)(MULT_SIZE-1) & MULT_83(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(3)(MULT_SIZE-1) & MULT_84(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(4)<=signed(MULT_83(4)(MULT_SIZE-1) & MULT_83(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(4)(MULT_SIZE-1) & MULT_84(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(5)<=signed(MULT_83(5)(MULT_SIZE-1) & MULT_83(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(5)(MULT_SIZE-1) & MULT_84(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(6)<=signed(MULT_83(6)(MULT_SIZE-1) & MULT_83(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(6)(MULT_SIZE-1) & MULT_84(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(7)<=signed(MULT_83(7)(MULT_SIZE-1) & MULT_83(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(7)(MULT_SIZE-1) & MULT_84(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(8)<=signed(MULT_83(8)(MULT_SIZE-1) & MULT_83(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(8)(MULT_SIZE-1) & MULT_84(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(9)<=signed(MULT_83(9)(MULT_SIZE-1) & MULT_83(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(9)(MULT_SIZE-1) & MULT_84(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));



                     EN_SUM_MULT_2<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_2 = '1' then
			------------------------------------STAGE-2--------------------------------------
			MULTS_2_1(0)<=signed(MULTS_1_1(0)(PERCISION) & MULTS_1_1(0)(PERCISION downto 1))+signed(MULTS_1_2(0)(PERCISION) & MULTS_1_2(0)(PERCISION downto 1));
			MULTS_2_1(1)<=signed(MULTS_1_1(1)(PERCISION) & MULTS_1_1(1)(PERCISION downto 1))+signed(MULTS_1_2(1)(PERCISION) & MULTS_1_2(1)(PERCISION downto 1));
			MULTS_2_1(2)<=signed(MULTS_1_1(2)(PERCISION) & MULTS_1_1(2)(PERCISION downto 1))+signed(MULTS_1_2(2)(PERCISION) & MULTS_1_2(2)(PERCISION downto 1));
			MULTS_2_1(3)<=signed(MULTS_1_1(3)(PERCISION) & MULTS_1_1(3)(PERCISION downto 1))+signed(MULTS_1_2(3)(PERCISION) & MULTS_1_2(3)(PERCISION downto 1));
			MULTS_2_1(4)<=signed(MULTS_1_1(4)(PERCISION) & MULTS_1_1(4)(PERCISION downto 1))+signed(MULTS_1_2(4)(PERCISION) & MULTS_1_2(4)(PERCISION downto 1));
			MULTS_2_1(5)<=signed(MULTS_1_1(5)(PERCISION) & MULTS_1_1(5)(PERCISION downto 1))+signed(MULTS_1_2(5)(PERCISION) & MULTS_1_2(5)(PERCISION downto 1));
			MULTS_2_1(6)<=signed(MULTS_1_1(6)(PERCISION) & MULTS_1_1(6)(PERCISION downto 1))+signed(MULTS_1_2(6)(PERCISION) & MULTS_1_2(6)(PERCISION downto 1));
			MULTS_2_1(7)<=signed(MULTS_1_1(7)(PERCISION) & MULTS_1_1(7)(PERCISION downto 1))+signed(MULTS_1_2(7)(PERCISION) & MULTS_1_2(7)(PERCISION downto 1));
			MULTS_2_1(8)<=signed(MULTS_1_1(8)(PERCISION) & MULTS_1_1(8)(PERCISION downto 1))+signed(MULTS_1_2(8)(PERCISION) & MULTS_1_2(8)(PERCISION downto 1));
			MULTS_2_1(9)<=signed(MULTS_1_1(9)(PERCISION) & MULTS_1_1(9)(PERCISION downto 1))+signed(MULTS_1_2(9)(PERCISION) & MULTS_1_2(9)(PERCISION downto 1));

			MULTS_2_2(0)<=signed(MULTS_1_3(0)(PERCISION) & MULTS_1_3(0)(PERCISION downto 1))+signed(MULTS_1_4(0)(PERCISION) & MULTS_1_4(0)(PERCISION downto 1));
			MULTS_2_2(1)<=signed(MULTS_1_3(1)(PERCISION) & MULTS_1_3(1)(PERCISION downto 1))+signed(MULTS_1_4(1)(PERCISION) & MULTS_1_4(1)(PERCISION downto 1));
			MULTS_2_2(2)<=signed(MULTS_1_3(2)(PERCISION) & MULTS_1_3(2)(PERCISION downto 1))+signed(MULTS_1_4(2)(PERCISION) & MULTS_1_4(2)(PERCISION downto 1));
			MULTS_2_2(3)<=signed(MULTS_1_3(3)(PERCISION) & MULTS_1_3(3)(PERCISION downto 1))+signed(MULTS_1_4(3)(PERCISION) & MULTS_1_4(3)(PERCISION downto 1));
			MULTS_2_2(4)<=signed(MULTS_1_3(4)(PERCISION) & MULTS_1_3(4)(PERCISION downto 1))+signed(MULTS_1_4(4)(PERCISION) & MULTS_1_4(4)(PERCISION downto 1));
			MULTS_2_2(5)<=signed(MULTS_1_3(5)(PERCISION) & MULTS_1_3(5)(PERCISION downto 1))+signed(MULTS_1_4(5)(PERCISION) & MULTS_1_4(5)(PERCISION downto 1));
			MULTS_2_2(6)<=signed(MULTS_1_3(6)(PERCISION) & MULTS_1_3(6)(PERCISION downto 1))+signed(MULTS_1_4(6)(PERCISION) & MULTS_1_4(6)(PERCISION downto 1));
			MULTS_2_2(7)<=signed(MULTS_1_3(7)(PERCISION) & MULTS_1_3(7)(PERCISION downto 1))+signed(MULTS_1_4(7)(PERCISION) & MULTS_1_4(7)(PERCISION downto 1));
			MULTS_2_2(8)<=signed(MULTS_1_3(8)(PERCISION) & MULTS_1_3(8)(PERCISION downto 1))+signed(MULTS_1_4(8)(PERCISION) & MULTS_1_4(8)(PERCISION downto 1));
			MULTS_2_2(9)<=signed(MULTS_1_3(9)(PERCISION) & MULTS_1_3(9)(PERCISION downto 1))+signed(MULTS_1_4(9)(PERCISION) & MULTS_1_4(9)(PERCISION downto 1));

			MULTS_2_3(0)<=signed(MULTS_1_5(0)(PERCISION) & MULTS_1_5(0)(PERCISION downto 1))+signed(MULTS_1_6(0)(PERCISION) & MULTS_1_6(0)(PERCISION downto 1));
			MULTS_2_3(1)<=signed(MULTS_1_5(1)(PERCISION) & MULTS_1_5(1)(PERCISION downto 1))+signed(MULTS_1_6(1)(PERCISION) & MULTS_1_6(1)(PERCISION downto 1));
			MULTS_2_3(2)<=signed(MULTS_1_5(2)(PERCISION) & MULTS_1_5(2)(PERCISION downto 1))+signed(MULTS_1_6(2)(PERCISION) & MULTS_1_6(2)(PERCISION downto 1));
			MULTS_2_3(3)<=signed(MULTS_1_5(3)(PERCISION) & MULTS_1_5(3)(PERCISION downto 1))+signed(MULTS_1_6(3)(PERCISION) & MULTS_1_6(3)(PERCISION downto 1));
			MULTS_2_3(4)<=signed(MULTS_1_5(4)(PERCISION) & MULTS_1_5(4)(PERCISION downto 1))+signed(MULTS_1_6(4)(PERCISION) & MULTS_1_6(4)(PERCISION downto 1));
			MULTS_2_3(5)<=signed(MULTS_1_5(5)(PERCISION) & MULTS_1_5(5)(PERCISION downto 1))+signed(MULTS_1_6(5)(PERCISION) & MULTS_1_6(5)(PERCISION downto 1));
			MULTS_2_3(6)<=signed(MULTS_1_5(6)(PERCISION) & MULTS_1_5(6)(PERCISION downto 1))+signed(MULTS_1_6(6)(PERCISION) & MULTS_1_6(6)(PERCISION downto 1));
			MULTS_2_3(7)<=signed(MULTS_1_5(7)(PERCISION) & MULTS_1_5(7)(PERCISION downto 1))+signed(MULTS_1_6(7)(PERCISION) & MULTS_1_6(7)(PERCISION downto 1));
			MULTS_2_3(8)<=signed(MULTS_1_5(8)(PERCISION) & MULTS_1_5(8)(PERCISION downto 1))+signed(MULTS_1_6(8)(PERCISION) & MULTS_1_6(8)(PERCISION downto 1));
			MULTS_2_3(9)<=signed(MULTS_1_5(9)(PERCISION) & MULTS_1_5(9)(PERCISION downto 1))+signed(MULTS_1_6(9)(PERCISION) & MULTS_1_6(9)(PERCISION downto 1));

			MULTS_2_4(0)<=signed(MULTS_1_7(0)(PERCISION) & MULTS_1_7(0)(PERCISION downto 1))+signed(MULTS_1_8(0)(PERCISION) & MULTS_1_8(0)(PERCISION downto 1));
			MULTS_2_4(1)<=signed(MULTS_1_7(1)(PERCISION) & MULTS_1_7(1)(PERCISION downto 1))+signed(MULTS_1_8(1)(PERCISION) & MULTS_1_8(1)(PERCISION downto 1));
			MULTS_2_4(2)<=signed(MULTS_1_7(2)(PERCISION) & MULTS_1_7(2)(PERCISION downto 1))+signed(MULTS_1_8(2)(PERCISION) & MULTS_1_8(2)(PERCISION downto 1));
			MULTS_2_4(3)<=signed(MULTS_1_7(3)(PERCISION) & MULTS_1_7(3)(PERCISION downto 1))+signed(MULTS_1_8(3)(PERCISION) & MULTS_1_8(3)(PERCISION downto 1));
			MULTS_2_4(4)<=signed(MULTS_1_7(4)(PERCISION) & MULTS_1_7(4)(PERCISION downto 1))+signed(MULTS_1_8(4)(PERCISION) & MULTS_1_8(4)(PERCISION downto 1));
			MULTS_2_4(5)<=signed(MULTS_1_7(5)(PERCISION) & MULTS_1_7(5)(PERCISION downto 1))+signed(MULTS_1_8(5)(PERCISION) & MULTS_1_8(5)(PERCISION downto 1));
			MULTS_2_4(6)<=signed(MULTS_1_7(6)(PERCISION) & MULTS_1_7(6)(PERCISION downto 1))+signed(MULTS_1_8(6)(PERCISION) & MULTS_1_8(6)(PERCISION downto 1));
			MULTS_2_4(7)<=signed(MULTS_1_7(7)(PERCISION) & MULTS_1_7(7)(PERCISION downto 1))+signed(MULTS_1_8(7)(PERCISION) & MULTS_1_8(7)(PERCISION downto 1));
			MULTS_2_4(8)<=signed(MULTS_1_7(8)(PERCISION) & MULTS_1_7(8)(PERCISION downto 1))+signed(MULTS_1_8(8)(PERCISION) & MULTS_1_8(8)(PERCISION downto 1));
			MULTS_2_4(9)<=signed(MULTS_1_7(9)(PERCISION) & MULTS_1_7(9)(PERCISION downto 1))+signed(MULTS_1_8(9)(PERCISION) & MULTS_1_8(9)(PERCISION downto 1));

			MULTS_2_5(0)<=signed(MULTS_1_9(0)(PERCISION) & MULTS_1_9(0)(PERCISION downto 1))+signed(MULTS_1_10(0)(PERCISION) & MULTS_1_10(0)(PERCISION downto 1));
			MULTS_2_5(1)<=signed(MULTS_1_9(1)(PERCISION) & MULTS_1_9(1)(PERCISION downto 1))+signed(MULTS_1_10(1)(PERCISION) & MULTS_1_10(1)(PERCISION downto 1));
			MULTS_2_5(2)<=signed(MULTS_1_9(2)(PERCISION) & MULTS_1_9(2)(PERCISION downto 1))+signed(MULTS_1_10(2)(PERCISION) & MULTS_1_10(2)(PERCISION downto 1));
			MULTS_2_5(3)<=signed(MULTS_1_9(3)(PERCISION) & MULTS_1_9(3)(PERCISION downto 1))+signed(MULTS_1_10(3)(PERCISION) & MULTS_1_10(3)(PERCISION downto 1));
			MULTS_2_5(4)<=signed(MULTS_1_9(4)(PERCISION) & MULTS_1_9(4)(PERCISION downto 1))+signed(MULTS_1_10(4)(PERCISION) & MULTS_1_10(4)(PERCISION downto 1));
			MULTS_2_5(5)<=signed(MULTS_1_9(5)(PERCISION) & MULTS_1_9(5)(PERCISION downto 1))+signed(MULTS_1_10(5)(PERCISION) & MULTS_1_10(5)(PERCISION downto 1));
			MULTS_2_5(6)<=signed(MULTS_1_9(6)(PERCISION) & MULTS_1_9(6)(PERCISION downto 1))+signed(MULTS_1_10(6)(PERCISION) & MULTS_1_10(6)(PERCISION downto 1));
			MULTS_2_5(7)<=signed(MULTS_1_9(7)(PERCISION) & MULTS_1_9(7)(PERCISION downto 1))+signed(MULTS_1_10(7)(PERCISION) & MULTS_1_10(7)(PERCISION downto 1));
			MULTS_2_5(8)<=signed(MULTS_1_9(8)(PERCISION) & MULTS_1_9(8)(PERCISION downto 1))+signed(MULTS_1_10(8)(PERCISION) & MULTS_1_10(8)(PERCISION downto 1));
			MULTS_2_5(9)<=signed(MULTS_1_9(9)(PERCISION) & MULTS_1_9(9)(PERCISION downto 1))+signed(MULTS_1_10(9)(PERCISION) & MULTS_1_10(9)(PERCISION downto 1));

			MULTS_2_6(0)<=signed(MULTS_1_11(0)(PERCISION) & MULTS_1_11(0)(PERCISION downto 1))+signed(MULTS_1_12(0)(PERCISION) & MULTS_1_12(0)(PERCISION downto 1));
			MULTS_2_6(1)<=signed(MULTS_1_11(1)(PERCISION) & MULTS_1_11(1)(PERCISION downto 1))+signed(MULTS_1_12(1)(PERCISION) & MULTS_1_12(1)(PERCISION downto 1));
			MULTS_2_6(2)<=signed(MULTS_1_11(2)(PERCISION) & MULTS_1_11(2)(PERCISION downto 1))+signed(MULTS_1_12(2)(PERCISION) & MULTS_1_12(2)(PERCISION downto 1));
			MULTS_2_6(3)<=signed(MULTS_1_11(3)(PERCISION) & MULTS_1_11(3)(PERCISION downto 1))+signed(MULTS_1_12(3)(PERCISION) & MULTS_1_12(3)(PERCISION downto 1));
			MULTS_2_6(4)<=signed(MULTS_1_11(4)(PERCISION) & MULTS_1_11(4)(PERCISION downto 1))+signed(MULTS_1_12(4)(PERCISION) & MULTS_1_12(4)(PERCISION downto 1));
			MULTS_2_6(5)<=signed(MULTS_1_11(5)(PERCISION) & MULTS_1_11(5)(PERCISION downto 1))+signed(MULTS_1_12(5)(PERCISION) & MULTS_1_12(5)(PERCISION downto 1));
			MULTS_2_6(6)<=signed(MULTS_1_11(6)(PERCISION) & MULTS_1_11(6)(PERCISION downto 1))+signed(MULTS_1_12(6)(PERCISION) & MULTS_1_12(6)(PERCISION downto 1));
			MULTS_2_6(7)<=signed(MULTS_1_11(7)(PERCISION) & MULTS_1_11(7)(PERCISION downto 1))+signed(MULTS_1_12(7)(PERCISION) & MULTS_1_12(7)(PERCISION downto 1));
			MULTS_2_6(8)<=signed(MULTS_1_11(8)(PERCISION) & MULTS_1_11(8)(PERCISION downto 1))+signed(MULTS_1_12(8)(PERCISION) & MULTS_1_12(8)(PERCISION downto 1));
			MULTS_2_6(9)<=signed(MULTS_1_11(9)(PERCISION) & MULTS_1_11(9)(PERCISION downto 1))+signed(MULTS_1_12(9)(PERCISION) & MULTS_1_12(9)(PERCISION downto 1));

			MULTS_2_7(0)<=signed(MULTS_1_13(0)(PERCISION) & MULTS_1_13(0)(PERCISION downto 1))+signed(MULTS_1_14(0)(PERCISION) & MULTS_1_14(0)(PERCISION downto 1));
			MULTS_2_7(1)<=signed(MULTS_1_13(1)(PERCISION) & MULTS_1_13(1)(PERCISION downto 1))+signed(MULTS_1_14(1)(PERCISION) & MULTS_1_14(1)(PERCISION downto 1));
			MULTS_2_7(2)<=signed(MULTS_1_13(2)(PERCISION) & MULTS_1_13(2)(PERCISION downto 1))+signed(MULTS_1_14(2)(PERCISION) & MULTS_1_14(2)(PERCISION downto 1));
			MULTS_2_7(3)<=signed(MULTS_1_13(3)(PERCISION) & MULTS_1_13(3)(PERCISION downto 1))+signed(MULTS_1_14(3)(PERCISION) & MULTS_1_14(3)(PERCISION downto 1));
			MULTS_2_7(4)<=signed(MULTS_1_13(4)(PERCISION) & MULTS_1_13(4)(PERCISION downto 1))+signed(MULTS_1_14(4)(PERCISION) & MULTS_1_14(4)(PERCISION downto 1));
			MULTS_2_7(5)<=signed(MULTS_1_13(5)(PERCISION) & MULTS_1_13(5)(PERCISION downto 1))+signed(MULTS_1_14(5)(PERCISION) & MULTS_1_14(5)(PERCISION downto 1));
			MULTS_2_7(6)<=signed(MULTS_1_13(6)(PERCISION) & MULTS_1_13(6)(PERCISION downto 1))+signed(MULTS_1_14(6)(PERCISION) & MULTS_1_14(6)(PERCISION downto 1));
			MULTS_2_7(7)<=signed(MULTS_1_13(7)(PERCISION) & MULTS_1_13(7)(PERCISION downto 1))+signed(MULTS_1_14(7)(PERCISION) & MULTS_1_14(7)(PERCISION downto 1));
			MULTS_2_7(8)<=signed(MULTS_1_13(8)(PERCISION) & MULTS_1_13(8)(PERCISION downto 1))+signed(MULTS_1_14(8)(PERCISION) & MULTS_1_14(8)(PERCISION downto 1));
			MULTS_2_7(9)<=signed(MULTS_1_13(9)(PERCISION) & MULTS_1_13(9)(PERCISION downto 1))+signed(MULTS_1_14(9)(PERCISION) & MULTS_1_14(9)(PERCISION downto 1));

			MULTS_2_8(0)<=signed(MULTS_1_15(0)(PERCISION) & MULTS_1_15(0)(PERCISION downto 1))+signed(MULTS_1_16(0)(PERCISION) & MULTS_1_16(0)(PERCISION downto 1));
			MULTS_2_8(1)<=signed(MULTS_1_15(1)(PERCISION) & MULTS_1_15(1)(PERCISION downto 1))+signed(MULTS_1_16(1)(PERCISION) & MULTS_1_16(1)(PERCISION downto 1));
			MULTS_2_8(2)<=signed(MULTS_1_15(2)(PERCISION) & MULTS_1_15(2)(PERCISION downto 1))+signed(MULTS_1_16(2)(PERCISION) & MULTS_1_16(2)(PERCISION downto 1));
			MULTS_2_8(3)<=signed(MULTS_1_15(3)(PERCISION) & MULTS_1_15(3)(PERCISION downto 1))+signed(MULTS_1_16(3)(PERCISION) & MULTS_1_16(3)(PERCISION downto 1));
			MULTS_2_8(4)<=signed(MULTS_1_15(4)(PERCISION) & MULTS_1_15(4)(PERCISION downto 1))+signed(MULTS_1_16(4)(PERCISION) & MULTS_1_16(4)(PERCISION downto 1));
			MULTS_2_8(5)<=signed(MULTS_1_15(5)(PERCISION) & MULTS_1_15(5)(PERCISION downto 1))+signed(MULTS_1_16(5)(PERCISION) & MULTS_1_16(5)(PERCISION downto 1));
			MULTS_2_8(6)<=signed(MULTS_1_15(6)(PERCISION) & MULTS_1_15(6)(PERCISION downto 1))+signed(MULTS_1_16(6)(PERCISION) & MULTS_1_16(6)(PERCISION downto 1));
			MULTS_2_8(7)<=signed(MULTS_1_15(7)(PERCISION) & MULTS_1_15(7)(PERCISION downto 1))+signed(MULTS_1_16(7)(PERCISION) & MULTS_1_16(7)(PERCISION downto 1));
			MULTS_2_8(8)<=signed(MULTS_1_15(8)(PERCISION) & MULTS_1_15(8)(PERCISION downto 1))+signed(MULTS_1_16(8)(PERCISION) & MULTS_1_16(8)(PERCISION downto 1));
			MULTS_2_8(9)<=signed(MULTS_1_15(9)(PERCISION) & MULTS_1_15(9)(PERCISION downto 1))+signed(MULTS_1_16(9)(PERCISION) & MULTS_1_16(9)(PERCISION downto 1));

			MULTS_2_9(0)<=signed(MULTS_1_17(0)(PERCISION) & MULTS_1_17(0)(PERCISION downto 1))+signed(MULTS_1_18(0)(PERCISION) & MULTS_1_18(0)(PERCISION downto 1));
			MULTS_2_9(1)<=signed(MULTS_1_17(1)(PERCISION) & MULTS_1_17(1)(PERCISION downto 1))+signed(MULTS_1_18(1)(PERCISION) & MULTS_1_18(1)(PERCISION downto 1));
			MULTS_2_9(2)<=signed(MULTS_1_17(2)(PERCISION) & MULTS_1_17(2)(PERCISION downto 1))+signed(MULTS_1_18(2)(PERCISION) & MULTS_1_18(2)(PERCISION downto 1));
			MULTS_2_9(3)<=signed(MULTS_1_17(3)(PERCISION) & MULTS_1_17(3)(PERCISION downto 1))+signed(MULTS_1_18(3)(PERCISION) & MULTS_1_18(3)(PERCISION downto 1));
			MULTS_2_9(4)<=signed(MULTS_1_17(4)(PERCISION) & MULTS_1_17(4)(PERCISION downto 1))+signed(MULTS_1_18(4)(PERCISION) & MULTS_1_18(4)(PERCISION downto 1));
			MULTS_2_9(5)<=signed(MULTS_1_17(5)(PERCISION) & MULTS_1_17(5)(PERCISION downto 1))+signed(MULTS_1_18(5)(PERCISION) & MULTS_1_18(5)(PERCISION downto 1));
			MULTS_2_9(6)<=signed(MULTS_1_17(6)(PERCISION) & MULTS_1_17(6)(PERCISION downto 1))+signed(MULTS_1_18(6)(PERCISION) & MULTS_1_18(6)(PERCISION downto 1));
			MULTS_2_9(7)<=signed(MULTS_1_17(7)(PERCISION) & MULTS_1_17(7)(PERCISION downto 1))+signed(MULTS_1_18(7)(PERCISION) & MULTS_1_18(7)(PERCISION downto 1));
			MULTS_2_9(8)<=signed(MULTS_1_17(8)(PERCISION) & MULTS_1_17(8)(PERCISION downto 1))+signed(MULTS_1_18(8)(PERCISION) & MULTS_1_18(8)(PERCISION downto 1));
			MULTS_2_9(9)<=signed(MULTS_1_17(9)(PERCISION) & MULTS_1_17(9)(PERCISION downto 1))+signed(MULTS_1_18(9)(PERCISION) & MULTS_1_18(9)(PERCISION downto 1));

			MULTS_2_10(0)<=signed(MULTS_1_19(0)(PERCISION) & MULTS_1_19(0)(PERCISION downto 1))+signed(MULTS_1_20(0)(PERCISION) & MULTS_1_20(0)(PERCISION downto 1));
			MULTS_2_10(1)<=signed(MULTS_1_19(1)(PERCISION) & MULTS_1_19(1)(PERCISION downto 1))+signed(MULTS_1_20(1)(PERCISION) & MULTS_1_20(1)(PERCISION downto 1));
			MULTS_2_10(2)<=signed(MULTS_1_19(2)(PERCISION) & MULTS_1_19(2)(PERCISION downto 1))+signed(MULTS_1_20(2)(PERCISION) & MULTS_1_20(2)(PERCISION downto 1));
			MULTS_2_10(3)<=signed(MULTS_1_19(3)(PERCISION) & MULTS_1_19(3)(PERCISION downto 1))+signed(MULTS_1_20(3)(PERCISION) & MULTS_1_20(3)(PERCISION downto 1));
			MULTS_2_10(4)<=signed(MULTS_1_19(4)(PERCISION) & MULTS_1_19(4)(PERCISION downto 1))+signed(MULTS_1_20(4)(PERCISION) & MULTS_1_20(4)(PERCISION downto 1));
			MULTS_2_10(5)<=signed(MULTS_1_19(5)(PERCISION) & MULTS_1_19(5)(PERCISION downto 1))+signed(MULTS_1_20(5)(PERCISION) & MULTS_1_20(5)(PERCISION downto 1));
			MULTS_2_10(6)<=signed(MULTS_1_19(6)(PERCISION) & MULTS_1_19(6)(PERCISION downto 1))+signed(MULTS_1_20(6)(PERCISION) & MULTS_1_20(6)(PERCISION downto 1));
			MULTS_2_10(7)<=signed(MULTS_1_19(7)(PERCISION) & MULTS_1_19(7)(PERCISION downto 1))+signed(MULTS_1_20(7)(PERCISION) & MULTS_1_20(7)(PERCISION downto 1));
			MULTS_2_10(8)<=signed(MULTS_1_19(8)(PERCISION) & MULTS_1_19(8)(PERCISION downto 1))+signed(MULTS_1_20(8)(PERCISION) & MULTS_1_20(8)(PERCISION downto 1));
			MULTS_2_10(9)<=signed(MULTS_1_19(9)(PERCISION) & MULTS_1_19(9)(PERCISION downto 1))+signed(MULTS_1_20(9)(PERCISION) & MULTS_1_20(9)(PERCISION downto 1));

			MULTS_2_11(0)<=signed(MULTS_1_21(0)(PERCISION) & MULTS_1_21(0)(PERCISION downto 1))+signed(MULTS_1_22(0)(PERCISION) & MULTS_1_22(0)(PERCISION downto 1));
			MULTS_2_11(1)<=signed(MULTS_1_21(1)(PERCISION) & MULTS_1_21(1)(PERCISION downto 1))+signed(MULTS_1_22(1)(PERCISION) & MULTS_1_22(1)(PERCISION downto 1));
			MULTS_2_11(2)<=signed(MULTS_1_21(2)(PERCISION) & MULTS_1_21(2)(PERCISION downto 1))+signed(MULTS_1_22(2)(PERCISION) & MULTS_1_22(2)(PERCISION downto 1));
			MULTS_2_11(3)<=signed(MULTS_1_21(3)(PERCISION) & MULTS_1_21(3)(PERCISION downto 1))+signed(MULTS_1_22(3)(PERCISION) & MULTS_1_22(3)(PERCISION downto 1));
			MULTS_2_11(4)<=signed(MULTS_1_21(4)(PERCISION) & MULTS_1_21(4)(PERCISION downto 1))+signed(MULTS_1_22(4)(PERCISION) & MULTS_1_22(4)(PERCISION downto 1));
			MULTS_2_11(5)<=signed(MULTS_1_21(5)(PERCISION) & MULTS_1_21(5)(PERCISION downto 1))+signed(MULTS_1_22(5)(PERCISION) & MULTS_1_22(5)(PERCISION downto 1));
			MULTS_2_11(6)<=signed(MULTS_1_21(6)(PERCISION) & MULTS_1_21(6)(PERCISION downto 1))+signed(MULTS_1_22(6)(PERCISION) & MULTS_1_22(6)(PERCISION downto 1));
			MULTS_2_11(7)<=signed(MULTS_1_21(7)(PERCISION) & MULTS_1_21(7)(PERCISION downto 1))+signed(MULTS_1_22(7)(PERCISION) & MULTS_1_22(7)(PERCISION downto 1));
			MULTS_2_11(8)<=signed(MULTS_1_21(8)(PERCISION) & MULTS_1_21(8)(PERCISION downto 1))+signed(MULTS_1_22(8)(PERCISION) & MULTS_1_22(8)(PERCISION downto 1));
			MULTS_2_11(9)<=signed(MULTS_1_21(9)(PERCISION) & MULTS_1_21(9)(PERCISION downto 1))+signed(MULTS_1_22(9)(PERCISION) & MULTS_1_22(9)(PERCISION downto 1));



                         EN_SUM_MULT_3<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_3 = '1' then
			------------------------------------STAGE-3--------------------------------------
			MULTS_3_1(0)<=signed(MULTS_2_1(0));
			MULTS_3_1(1)<=signed(MULTS_2_1(1));
			MULTS_3_1(2)<=signed(MULTS_2_1(2));
			MULTS_3_1(3)<=signed(MULTS_2_1(3));
			MULTS_3_1(4)<=signed(MULTS_2_1(4));
			MULTS_3_1(5)<=signed(MULTS_2_1(5));
			MULTS_3_1(6)<=signed(MULTS_2_1(6));
			MULTS_3_1(7)<=signed(MULTS_2_1(7));
			MULTS_3_1(8)<=signed(MULTS_2_1(8));
			MULTS_3_1(9)<=signed(MULTS_2_1(9));

			MULTS_3_2(0)<=signed(MULTS_2_2(0)(PERCISION) & MULTS_2_2(0)(PERCISION downto 1))+signed(MULTS_2_3(0)(PERCISION) & MULTS_2_3(0)(PERCISION downto 1));
			MULTS_3_2(1)<=signed(MULTS_2_2(1)(PERCISION) & MULTS_2_2(1)(PERCISION downto 1))+signed(MULTS_2_3(1)(PERCISION) & MULTS_2_3(1)(PERCISION downto 1));
			MULTS_3_2(2)<=signed(MULTS_2_2(2)(PERCISION) & MULTS_2_2(2)(PERCISION downto 1))+signed(MULTS_2_3(2)(PERCISION) & MULTS_2_3(2)(PERCISION downto 1));
			MULTS_3_2(3)<=signed(MULTS_2_2(3)(PERCISION) & MULTS_2_2(3)(PERCISION downto 1))+signed(MULTS_2_3(3)(PERCISION) & MULTS_2_3(3)(PERCISION downto 1));
			MULTS_3_2(4)<=signed(MULTS_2_2(4)(PERCISION) & MULTS_2_2(4)(PERCISION downto 1))+signed(MULTS_2_3(4)(PERCISION) & MULTS_2_3(4)(PERCISION downto 1));
			MULTS_3_2(5)<=signed(MULTS_2_2(5)(PERCISION) & MULTS_2_2(5)(PERCISION downto 1))+signed(MULTS_2_3(5)(PERCISION) & MULTS_2_3(5)(PERCISION downto 1));
			MULTS_3_2(6)<=signed(MULTS_2_2(6)(PERCISION) & MULTS_2_2(6)(PERCISION downto 1))+signed(MULTS_2_3(6)(PERCISION) & MULTS_2_3(6)(PERCISION downto 1));
			MULTS_3_2(7)<=signed(MULTS_2_2(7)(PERCISION) & MULTS_2_2(7)(PERCISION downto 1))+signed(MULTS_2_3(7)(PERCISION) & MULTS_2_3(7)(PERCISION downto 1));
			MULTS_3_2(8)<=signed(MULTS_2_2(8)(PERCISION) & MULTS_2_2(8)(PERCISION downto 1))+signed(MULTS_2_3(8)(PERCISION) & MULTS_2_3(8)(PERCISION downto 1));
			MULTS_3_2(9)<=signed(MULTS_2_2(9)(PERCISION) & MULTS_2_2(9)(PERCISION downto 1))+signed(MULTS_2_3(9)(PERCISION) & MULTS_2_3(9)(PERCISION downto 1));

			MULTS_3_3(0)<=signed(MULTS_2_4(0)(PERCISION) & MULTS_2_4(0)(PERCISION downto 1))+signed(MULTS_2_5(0)(PERCISION) & MULTS_2_5(0)(PERCISION downto 1));
			MULTS_3_3(1)<=signed(MULTS_2_4(1)(PERCISION) & MULTS_2_4(1)(PERCISION downto 1))+signed(MULTS_2_5(1)(PERCISION) & MULTS_2_5(1)(PERCISION downto 1));
			MULTS_3_3(2)<=signed(MULTS_2_4(2)(PERCISION) & MULTS_2_4(2)(PERCISION downto 1))+signed(MULTS_2_5(2)(PERCISION) & MULTS_2_5(2)(PERCISION downto 1));
			MULTS_3_3(3)<=signed(MULTS_2_4(3)(PERCISION) & MULTS_2_4(3)(PERCISION downto 1))+signed(MULTS_2_5(3)(PERCISION) & MULTS_2_5(3)(PERCISION downto 1));
			MULTS_3_3(4)<=signed(MULTS_2_4(4)(PERCISION) & MULTS_2_4(4)(PERCISION downto 1))+signed(MULTS_2_5(4)(PERCISION) & MULTS_2_5(4)(PERCISION downto 1));
			MULTS_3_3(5)<=signed(MULTS_2_4(5)(PERCISION) & MULTS_2_4(5)(PERCISION downto 1))+signed(MULTS_2_5(5)(PERCISION) & MULTS_2_5(5)(PERCISION downto 1));
			MULTS_3_3(6)<=signed(MULTS_2_4(6)(PERCISION) & MULTS_2_4(6)(PERCISION downto 1))+signed(MULTS_2_5(6)(PERCISION) & MULTS_2_5(6)(PERCISION downto 1));
			MULTS_3_3(7)<=signed(MULTS_2_4(7)(PERCISION) & MULTS_2_4(7)(PERCISION downto 1))+signed(MULTS_2_5(7)(PERCISION) & MULTS_2_5(7)(PERCISION downto 1));
			MULTS_3_3(8)<=signed(MULTS_2_4(8)(PERCISION) & MULTS_2_4(8)(PERCISION downto 1))+signed(MULTS_2_5(8)(PERCISION) & MULTS_2_5(8)(PERCISION downto 1));
			MULTS_3_3(9)<=signed(MULTS_2_4(9)(PERCISION) & MULTS_2_4(9)(PERCISION downto 1))+signed(MULTS_2_5(9)(PERCISION) & MULTS_2_5(9)(PERCISION downto 1));

			MULTS_3_4(0)<=signed(MULTS_2_6(0)(PERCISION) & MULTS_2_6(0)(PERCISION downto 1))+signed(MULTS_2_7(0)(PERCISION) & MULTS_2_7(0)(PERCISION downto 1));
			MULTS_3_4(1)<=signed(MULTS_2_6(1)(PERCISION) & MULTS_2_6(1)(PERCISION downto 1))+signed(MULTS_2_7(1)(PERCISION) & MULTS_2_7(1)(PERCISION downto 1));
			MULTS_3_4(2)<=signed(MULTS_2_6(2)(PERCISION) & MULTS_2_6(2)(PERCISION downto 1))+signed(MULTS_2_7(2)(PERCISION) & MULTS_2_7(2)(PERCISION downto 1));
			MULTS_3_4(3)<=signed(MULTS_2_6(3)(PERCISION) & MULTS_2_6(3)(PERCISION downto 1))+signed(MULTS_2_7(3)(PERCISION) & MULTS_2_7(3)(PERCISION downto 1));
			MULTS_3_4(4)<=signed(MULTS_2_6(4)(PERCISION) & MULTS_2_6(4)(PERCISION downto 1))+signed(MULTS_2_7(4)(PERCISION) & MULTS_2_7(4)(PERCISION downto 1));
			MULTS_3_4(5)<=signed(MULTS_2_6(5)(PERCISION) & MULTS_2_6(5)(PERCISION downto 1))+signed(MULTS_2_7(5)(PERCISION) & MULTS_2_7(5)(PERCISION downto 1));
			MULTS_3_4(6)<=signed(MULTS_2_6(6)(PERCISION) & MULTS_2_6(6)(PERCISION downto 1))+signed(MULTS_2_7(6)(PERCISION) & MULTS_2_7(6)(PERCISION downto 1));
			MULTS_3_4(7)<=signed(MULTS_2_6(7)(PERCISION) & MULTS_2_6(7)(PERCISION downto 1))+signed(MULTS_2_7(7)(PERCISION) & MULTS_2_7(7)(PERCISION downto 1));
			MULTS_3_4(8)<=signed(MULTS_2_6(8)(PERCISION) & MULTS_2_6(8)(PERCISION downto 1))+signed(MULTS_2_7(8)(PERCISION) & MULTS_2_7(8)(PERCISION downto 1));
			MULTS_3_4(9)<=signed(MULTS_2_6(9)(PERCISION) & MULTS_2_6(9)(PERCISION downto 1))+signed(MULTS_2_7(9)(PERCISION) & MULTS_2_7(9)(PERCISION downto 1));

			MULTS_3_5(0)<=signed(MULTS_2_8(0)(PERCISION) & MULTS_2_8(0)(PERCISION downto 1))+signed(MULTS_2_9(0)(PERCISION) & MULTS_2_9(0)(PERCISION downto 1));
			MULTS_3_5(1)<=signed(MULTS_2_8(1)(PERCISION) & MULTS_2_8(1)(PERCISION downto 1))+signed(MULTS_2_9(1)(PERCISION) & MULTS_2_9(1)(PERCISION downto 1));
			MULTS_3_5(2)<=signed(MULTS_2_8(2)(PERCISION) & MULTS_2_8(2)(PERCISION downto 1))+signed(MULTS_2_9(2)(PERCISION) & MULTS_2_9(2)(PERCISION downto 1));
			MULTS_3_5(3)<=signed(MULTS_2_8(3)(PERCISION) & MULTS_2_8(3)(PERCISION downto 1))+signed(MULTS_2_9(3)(PERCISION) & MULTS_2_9(3)(PERCISION downto 1));
			MULTS_3_5(4)<=signed(MULTS_2_8(4)(PERCISION) & MULTS_2_8(4)(PERCISION downto 1))+signed(MULTS_2_9(4)(PERCISION) & MULTS_2_9(4)(PERCISION downto 1));
			MULTS_3_5(5)<=signed(MULTS_2_8(5)(PERCISION) & MULTS_2_8(5)(PERCISION downto 1))+signed(MULTS_2_9(5)(PERCISION) & MULTS_2_9(5)(PERCISION downto 1));
			MULTS_3_5(6)<=signed(MULTS_2_8(6)(PERCISION) & MULTS_2_8(6)(PERCISION downto 1))+signed(MULTS_2_9(6)(PERCISION) & MULTS_2_9(6)(PERCISION downto 1));
			MULTS_3_5(7)<=signed(MULTS_2_8(7)(PERCISION) & MULTS_2_8(7)(PERCISION downto 1))+signed(MULTS_2_9(7)(PERCISION) & MULTS_2_9(7)(PERCISION downto 1));
			MULTS_3_5(8)<=signed(MULTS_2_8(8)(PERCISION) & MULTS_2_8(8)(PERCISION downto 1))+signed(MULTS_2_9(8)(PERCISION) & MULTS_2_9(8)(PERCISION downto 1));
			MULTS_3_5(9)<=signed(MULTS_2_8(9)(PERCISION) & MULTS_2_8(9)(PERCISION downto 1))+signed(MULTS_2_9(9)(PERCISION) & MULTS_2_9(9)(PERCISION downto 1));

			MULTS_3_6(0)<=signed(MULTS_2_10(0)(PERCISION) & MULTS_2_10(0)(PERCISION downto 1))+signed(MULTS_2_11(0)(PERCISION) & MULTS_2_11(0)(PERCISION downto 1));
			MULTS_3_6(1)<=signed(MULTS_2_10(1)(PERCISION) & MULTS_2_10(1)(PERCISION downto 1))+signed(MULTS_2_11(1)(PERCISION) & MULTS_2_11(1)(PERCISION downto 1));
			MULTS_3_6(2)<=signed(MULTS_2_10(2)(PERCISION) & MULTS_2_10(2)(PERCISION downto 1))+signed(MULTS_2_11(2)(PERCISION) & MULTS_2_11(2)(PERCISION downto 1));
			MULTS_3_6(3)<=signed(MULTS_2_10(3)(PERCISION) & MULTS_2_10(3)(PERCISION downto 1))+signed(MULTS_2_11(3)(PERCISION) & MULTS_2_11(3)(PERCISION downto 1));
			MULTS_3_6(4)<=signed(MULTS_2_10(4)(PERCISION) & MULTS_2_10(4)(PERCISION downto 1))+signed(MULTS_2_11(4)(PERCISION) & MULTS_2_11(4)(PERCISION downto 1));
			MULTS_3_6(5)<=signed(MULTS_2_10(5)(PERCISION) & MULTS_2_10(5)(PERCISION downto 1))+signed(MULTS_2_11(5)(PERCISION) & MULTS_2_11(5)(PERCISION downto 1));
			MULTS_3_6(6)<=signed(MULTS_2_10(6)(PERCISION) & MULTS_2_10(6)(PERCISION downto 1))+signed(MULTS_2_11(6)(PERCISION) & MULTS_2_11(6)(PERCISION downto 1));
			MULTS_3_6(7)<=signed(MULTS_2_10(7)(PERCISION) & MULTS_2_10(7)(PERCISION downto 1))+signed(MULTS_2_11(7)(PERCISION) & MULTS_2_11(7)(PERCISION downto 1));
			MULTS_3_6(8)<=signed(MULTS_2_10(8)(PERCISION) & MULTS_2_10(8)(PERCISION downto 1))+signed(MULTS_2_11(8)(PERCISION) & MULTS_2_11(8)(PERCISION downto 1));
			MULTS_3_6(9)<=signed(MULTS_2_10(9)(PERCISION) & MULTS_2_10(9)(PERCISION downto 1))+signed(MULTS_2_11(9)(PERCISION) & MULTS_2_11(9)(PERCISION downto 1));



                         EN_SUM_MULT_4<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_4 = '1' then
			------------------------------------STAGE-4--------------------------------------
			MULTS_4_1(0)<=signed(MULTS_3_1(0));
			MULTS_4_1(1)<=signed(MULTS_3_1(1));
			MULTS_4_1(2)<=signed(MULTS_3_1(2));
			MULTS_4_1(3)<=signed(MULTS_3_1(3));
			MULTS_4_1(4)<=signed(MULTS_3_1(4));
			MULTS_4_1(5)<=signed(MULTS_3_1(5));
			MULTS_4_1(6)<=signed(MULTS_3_1(6));
			MULTS_4_1(7)<=signed(MULTS_3_1(7));
			MULTS_4_1(8)<=signed(MULTS_3_1(8));
			MULTS_4_1(9)<=signed(MULTS_3_1(9));

			MULTS_4_2(0)<=signed(MULTS_3_2(0)(PERCISION) & MULTS_3_2(0)(PERCISION downto 1))+signed(MULTS_3_3(0)(PERCISION) & MULTS_3_3(0)(PERCISION downto 1));
			MULTS_4_2(1)<=signed(MULTS_3_2(1)(PERCISION) & MULTS_3_2(1)(PERCISION downto 1))+signed(MULTS_3_3(1)(PERCISION) & MULTS_3_3(1)(PERCISION downto 1));
			MULTS_4_2(2)<=signed(MULTS_3_2(2)(PERCISION) & MULTS_3_2(2)(PERCISION downto 1))+signed(MULTS_3_3(2)(PERCISION) & MULTS_3_3(2)(PERCISION downto 1));
			MULTS_4_2(3)<=signed(MULTS_3_2(3)(PERCISION) & MULTS_3_2(3)(PERCISION downto 1))+signed(MULTS_3_3(3)(PERCISION) & MULTS_3_3(3)(PERCISION downto 1));
			MULTS_4_2(4)<=signed(MULTS_3_2(4)(PERCISION) & MULTS_3_2(4)(PERCISION downto 1))+signed(MULTS_3_3(4)(PERCISION) & MULTS_3_3(4)(PERCISION downto 1));
			MULTS_4_2(5)<=signed(MULTS_3_2(5)(PERCISION) & MULTS_3_2(5)(PERCISION downto 1))+signed(MULTS_3_3(5)(PERCISION) & MULTS_3_3(5)(PERCISION downto 1));
			MULTS_4_2(6)<=signed(MULTS_3_2(6)(PERCISION) & MULTS_3_2(6)(PERCISION downto 1))+signed(MULTS_3_3(6)(PERCISION) & MULTS_3_3(6)(PERCISION downto 1));
			MULTS_4_2(7)<=signed(MULTS_3_2(7)(PERCISION) & MULTS_3_2(7)(PERCISION downto 1))+signed(MULTS_3_3(7)(PERCISION) & MULTS_3_3(7)(PERCISION downto 1));
			MULTS_4_2(8)<=signed(MULTS_3_2(8)(PERCISION) & MULTS_3_2(8)(PERCISION downto 1))+signed(MULTS_3_3(8)(PERCISION) & MULTS_3_3(8)(PERCISION downto 1));
			MULTS_4_2(9)<=signed(MULTS_3_2(9)(PERCISION) & MULTS_3_2(9)(PERCISION downto 1))+signed(MULTS_3_3(9)(PERCISION) & MULTS_3_3(9)(PERCISION downto 1));

			MULTS_4_3(0)<=signed(MULTS_3_4(0)(PERCISION) & MULTS_3_4(0)(PERCISION downto 1))+signed(MULTS_3_5(0)(PERCISION) & MULTS_3_5(0)(PERCISION downto 1));
			MULTS_4_3(1)<=signed(MULTS_3_4(1)(PERCISION) & MULTS_3_4(1)(PERCISION downto 1))+signed(MULTS_3_5(1)(PERCISION) & MULTS_3_5(1)(PERCISION downto 1));
			MULTS_4_3(2)<=signed(MULTS_3_4(2)(PERCISION) & MULTS_3_4(2)(PERCISION downto 1))+signed(MULTS_3_5(2)(PERCISION) & MULTS_3_5(2)(PERCISION downto 1));
			MULTS_4_3(3)<=signed(MULTS_3_4(3)(PERCISION) & MULTS_3_4(3)(PERCISION downto 1))+signed(MULTS_3_5(3)(PERCISION) & MULTS_3_5(3)(PERCISION downto 1));
			MULTS_4_3(4)<=signed(MULTS_3_4(4)(PERCISION) & MULTS_3_4(4)(PERCISION downto 1))+signed(MULTS_3_5(4)(PERCISION) & MULTS_3_5(4)(PERCISION downto 1));
			MULTS_4_3(5)<=signed(MULTS_3_4(5)(PERCISION) & MULTS_3_4(5)(PERCISION downto 1))+signed(MULTS_3_5(5)(PERCISION) & MULTS_3_5(5)(PERCISION downto 1));
			MULTS_4_3(6)<=signed(MULTS_3_4(6)(PERCISION) & MULTS_3_4(6)(PERCISION downto 1))+signed(MULTS_3_5(6)(PERCISION) & MULTS_3_5(6)(PERCISION downto 1));
			MULTS_4_3(7)<=signed(MULTS_3_4(7)(PERCISION) & MULTS_3_4(7)(PERCISION downto 1))+signed(MULTS_3_5(7)(PERCISION) & MULTS_3_5(7)(PERCISION downto 1));
			MULTS_4_3(8)<=signed(MULTS_3_4(8)(PERCISION) & MULTS_3_4(8)(PERCISION downto 1))+signed(MULTS_3_5(8)(PERCISION) & MULTS_3_5(8)(PERCISION downto 1));
			MULTS_4_3(9)<=signed(MULTS_3_4(9)(PERCISION) & MULTS_3_4(9)(PERCISION downto 1))+signed(MULTS_3_5(9)(PERCISION) & MULTS_3_5(9)(PERCISION downto 1));

			MULTS_4_4(0)<=signed(MULTS_3_6(0)(PERCISION) & MULTS_3_6(0)(PERCISION downto 1))+signed(MULTS_3_7(0)(PERCISION) & MULTS_3_7(0)(PERCISION downto 1));
			MULTS_4_4(1)<=signed(MULTS_3_6(1)(PERCISION) & MULTS_3_6(1)(PERCISION downto 1))+signed(MULTS_3_7(1)(PERCISION) & MULTS_3_7(1)(PERCISION downto 1));
			MULTS_4_4(2)<=signed(MULTS_3_6(2)(PERCISION) & MULTS_3_6(2)(PERCISION downto 1))+signed(MULTS_3_7(2)(PERCISION) & MULTS_3_7(2)(PERCISION downto 1));
			MULTS_4_4(3)<=signed(MULTS_3_6(3)(PERCISION) & MULTS_3_6(3)(PERCISION downto 1))+signed(MULTS_3_7(3)(PERCISION) & MULTS_3_7(3)(PERCISION downto 1));
			MULTS_4_4(4)<=signed(MULTS_3_6(4)(PERCISION) & MULTS_3_6(4)(PERCISION downto 1))+signed(MULTS_3_7(4)(PERCISION) & MULTS_3_7(4)(PERCISION downto 1));
			MULTS_4_4(5)<=signed(MULTS_3_6(5)(PERCISION) & MULTS_3_6(5)(PERCISION downto 1))+signed(MULTS_3_7(5)(PERCISION) & MULTS_3_7(5)(PERCISION downto 1));
			MULTS_4_4(6)<=signed(MULTS_3_6(6)(PERCISION) & MULTS_3_6(6)(PERCISION downto 1))+signed(MULTS_3_7(6)(PERCISION) & MULTS_3_7(6)(PERCISION downto 1));
			MULTS_4_4(7)<=signed(MULTS_3_6(7)(PERCISION) & MULTS_3_6(7)(PERCISION downto 1))+signed(MULTS_3_7(7)(PERCISION) & MULTS_3_7(7)(PERCISION downto 1));
			MULTS_4_4(8)<=signed(MULTS_3_6(8)(PERCISION) & MULTS_3_6(8)(PERCISION downto 1))+signed(MULTS_3_7(8)(PERCISION) & MULTS_3_7(8)(PERCISION downto 1));
			MULTS_4_4(9)<=signed(MULTS_3_6(9)(PERCISION) & MULTS_3_6(9)(PERCISION downto 1))+signed(MULTS_3_7(9)(PERCISION) & MULTS_3_7(9)(PERCISION downto 1));



                         EN_SUM_MULT_5<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_5 = '1' then
			------------------------------------STAGE-5--------------------------------------
			MULTS_5_1(0)<=signed(MULTS_4_1(0)(PERCISION) & MULTS_4_1(0)(PERCISION downto 1))+signed(MULTS_4_2(0)(PERCISION) & MULTS_4_2(0)(PERCISION downto 1));
			MULTS_5_1(1)<=signed(MULTS_4_1(1)(PERCISION) & MULTS_4_1(1)(PERCISION downto 1))+signed(MULTS_4_2(1)(PERCISION) & MULTS_4_2(1)(PERCISION downto 1));
			MULTS_5_1(2)<=signed(MULTS_4_1(2)(PERCISION) & MULTS_4_1(2)(PERCISION downto 1))+signed(MULTS_4_2(2)(PERCISION) & MULTS_4_2(2)(PERCISION downto 1));
			MULTS_5_1(3)<=signed(MULTS_4_1(3)(PERCISION) & MULTS_4_1(3)(PERCISION downto 1))+signed(MULTS_4_2(3)(PERCISION) & MULTS_4_2(3)(PERCISION downto 1));
			MULTS_5_1(4)<=signed(MULTS_4_1(4)(PERCISION) & MULTS_4_1(4)(PERCISION downto 1))+signed(MULTS_4_2(4)(PERCISION) & MULTS_4_2(4)(PERCISION downto 1));
			MULTS_5_1(5)<=signed(MULTS_4_1(5)(PERCISION) & MULTS_4_1(5)(PERCISION downto 1))+signed(MULTS_4_2(5)(PERCISION) & MULTS_4_2(5)(PERCISION downto 1));
			MULTS_5_1(6)<=signed(MULTS_4_1(6)(PERCISION) & MULTS_4_1(6)(PERCISION downto 1))+signed(MULTS_4_2(6)(PERCISION) & MULTS_4_2(6)(PERCISION downto 1));
			MULTS_5_1(7)<=signed(MULTS_4_1(7)(PERCISION) & MULTS_4_1(7)(PERCISION downto 1))+signed(MULTS_4_2(7)(PERCISION) & MULTS_4_2(7)(PERCISION downto 1));
			MULTS_5_1(8)<=signed(MULTS_4_1(8)(PERCISION) & MULTS_4_1(8)(PERCISION downto 1))+signed(MULTS_4_2(8)(PERCISION) & MULTS_4_2(8)(PERCISION downto 1));
			MULTS_5_1(9)<=signed(MULTS_4_1(9)(PERCISION) & MULTS_4_1(9)(PERCISION downto 1))+signed(MULTS_4_2(9)(PERCISION) & MULTS_4_2(9)(PERCISION downto 1));

			MULTS_5_2(0)<=signed(MULTS_4_3(0)(PERCISION) & MULTS_4_3(0)(PERCISION downto 1))+signed(MULTS_4_4(0)(PERCISION) & MULTS_4_4(0)(PERCISION downto 1));
			MULTS_5_2(1)<=signed(MULTS_4_3(1)(PERCISION) & MULTS_4_3(1)(PERCISION downto 1))+signed(MULTS_4_4(1)(PERCISION) & MULTS_4_4(1)(PERCISION downto 1));
			MULTS_5_2(2)<=signed(MULTS_4_3(2)(PERCISION) & MULTS_4_3(2)(PERCISION downto 1))+signed(MULTS_4_4(2)(PERCISION) & MULTS_4_4(2)(PERCISION downto 1));
			MULTS_5_2(3)<=signed(MULTS_4_3(3)(PERCISION) & MULTS_4_3(3)(PERCISION downto 1))+signed(MULTS_4_4(3)(PERCISION) & MULTS_4_4(3)(PERCISION downto 1));
			MULTS_5_2(4)<=signed(MULTS_4_3(4)(PERCISION) & MULTS_4_3(4)(PERCISION downto 1))+signed(MULTS_4_4(4)(PERCISION) & MULTS_4_4(4)(PERCISION downto 1));
			MULTS_5_2(5)<=signed(MULTS_4_3(5)(PERCISION) & MULTS_4_3(5)(PERCISION downto 1))+signed(MULTS_4_4(5)(PERCISION) & MULTS_4_4(5)(PERCISION downto 1));
			MULTS_5_2(6)<=signed(MULTS_4_3(6)(PERCISION) & MULTS_4_3(6)(PERCISION downto 1))+signed(MULTS_4_4(6)(PERCISION) & MULTS_4_4(6)(PERCISION downto 1));
			MULTS_5_2(7)<=signed(MULTS_4_3(7)(PERCISION) & MULTS_4_3(7)(PERCISION downto 1))+signed(MULTS_4_4(7)(PERCISION) & MULTS_4_4(7)(PERCISION downto 1));
			MULTS_5_2(8)<=signed(MULTS_4_3(8)(PERCISION) & MULTS_4_3(8)(PERCISION downto 1))+signed(MULTS_4_4(8)(PERCISION) & MULTS_4_4(8)(PERCISION downto 1));
			MULTS_5_2(9)<=signed(MULTS_4_3(9)(PERCISION) & MULTS_4_3(9)(PERCISION downto 1))+signed(MULTS_4_4(9)(PERCISION) & MULTS_4_4(9)(PERCISION downto 1));



                         EN_SUM_MULT_6<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_6 = '1' then
			------------------------------------STAGE-6--------------------------------------
			MULTS_6_1(0)<=signed(MULTS_5_1(0));
			MULTS_6_1(1)<=signed(MULTS_5_1(1));
			MULTS_6_1(2)<=signed(MULTS_5_1(2));
			MULTS_6_1(3)<=signed(MULTS_5_1(3));
			MULTS_6_1(4)<=signed(MULTS_5_1(4));
			MULTS_6_1(5)<=signed(MULTS_5_1(5));
			MULTS_6_1(6)<=signed(MULTS_5_1(6));
			MULTS_6_1(7)<=signed(MULTS_5_1(7));
			MULTS_6_1(8)<=signed(MULTS_5_1(8));
			MULTS_6_1(9)<=signed(MULTS_5_1(9));

			MULTS_6_2(0)<=signed(MULTS_5_2(0)(PERCISION) & MULTS_5_2(0)(PERCISION downto 1))+signed(MULTS_5_3(0)(PERCISION) & MULTS_5_3(0)(PERCISION downto 1));
			MULTS_6_2(1)<=signed(MULTS_5_2(1)(PERCISION) & MULTS_5_2(1)(PERCISION downto 1))+signed(MULTS_5_3(1)(PERCISION) & MULTS_5_3(1)(PERCISION downto 1));
			MULTS_6_2(2)<=signed(MULTS_5_2(2)(PERCISION) & MULTS_5_2(2)(PERCISION downto 1))+signed(MULTS_5_3(2)(PERCISION) & MULTS_5_3(2)(PERCISION downto 1));
			MULTS_6_2(3)<=signed(MULTS_5_2(3)(PERCISION) & MULTS_5_2(3)(PERCISION downto 1))+signed(MULTS_5_3(3)(PERCISION) & MULTS_5_3(3)(PERCISION downto 1));
			MULTS_6_2(4)<=signed(MULTS_5_2(4)(PERCISION) & MULTS_5_2(4)(PERCISION downto 1))+signed(MULTS_5_3(4)(PERCISION) & MULTS_5_3(4)(PERCISION downto 1));
			MULTS_6_2(5)<=signed(MULTS_5_2(5)(PERCISION) & MULTS_5_2(5)(PERCISION downto 1))+signed(MULTS_5_3(5)(PERCISION) & MULTS_5_3(5)(PERCISION downto 1));
			MULTS_6_2(6)<=signed(MULTS_5_2(6)(PERCISION) & MULTS_5_2(6)(PERCISION downto 1))+signed(MULTS_5_3(6)(PERCISION) & MULTS_5_3(6)(PERCISION downto 1));
			MULTS_6_2(7)<=signed(MULTS_5_2(7)(PERCISION) & MULTS_5_2(7)(PERCISION downto 1))+signed(MULTS_5_3(7)(PERCISION) & MULTS_5_3(7)(PERCISION downto 1));
			MULTS_6_2(8)<=signed(MULTS_5_2(8)(PERCISION) & MULTS_5_2(8)(PERCISION downto 1))+signed(MULTS_5_3(8)(PERCISION) & MULTS_5_3(8)(PERCISION downto 1));
			MULTS_6_2(9)<=signed(MULTS_5_2(9)(PERCISION) & MULTS_5_2(9)(PERCISION downto 1))+signed(MULTS_5_3(9)(PERCISION) & MULTS_5_3(9)(PERCISION downto 1));



                         EN_SUM_MULT_7<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_7 = '1' then
			------------------------------------STAGE-7--------------------------------------
			MULTS_7_1(0)<=signed(MULTS_6_1(0)(PERCISION) & MULTS_6_1(0)(PERCISION downto 1))+signed(MULTS_6_2(0)(PERCISION) & MULTS_6_2(0)(PERCISION downto 1));
			MULTS_7_1(1)<=signed(MULTS_6_1(1)(PERCISION) & MULTS_6_1(1)(PERCISION downto 1))+signed(MULTS_6_2(1)(PERCISION) & MULTS_6_2(1)(PERCISION downto 1));
			MULTS_7_1(2)<=signed(MULTS_6_1(2)(PERCISION) & MULTS_6_1(2)(PERCISION downto 1))+signed(MULTS_6_2(2)(PERCISION) & MULTS_6_2(2)(PERCISION downto 1));
			MULTS_7_1(3)<=signed(MULTS_6_1(3)(PERCISION) & MULTS_6_1(3)(PERCISION downto 1))+signed(MULTS_6_2(3)(PERCISION) & MULTS_6_2(3)(PERCISION downto 1));
			MULTS_7_1(4)<=signed(MULTS_6_1(4)(PERCISION) & MULTS_6_1(4)(PERCISION downto 1))+signed(MULTS_6_2(4)(PERCISION) & MULTS_6_2(4)(PERCISION downto 1));
			MULTS_7_1(5)<=signed(MULTS_6_1(5)(PERCISION) & MULTS_6_1(5)(PERCISION downto 1))+signed(MULTS_6_2(5)(PERCISION) & MULTS_6_2(5)(PERCISION downto 1));
			MULTS_7_1(6)<=signed(MULTS_6_1(6)(PERCISION) & MULTS_6_1(6)(PERCISION downto 1))+signed(MULTS_6_2(6)(PERCISION) & MULTS_6_2(6)(PERCISION downto 1));
			MULTS_7_1(7)<=signed(MULTS_6_1(7)(PERCISION) & MULTS_6_1(7)(PERCISION downto 1))+signed(MULTS_6_2(7)(PERCISION) & MULTS_6_2(7)(PERCISION downto 1));
			MULTS_7_1(8)<=signed(MULTS_6_1(8)(PERCISION) & MULTS_6_1(8)(PERCISION downto 1))+signed(MULTS_6_2(8)(PERCISION) & MULTS_6_2(8)(PERCISION downto 1));
			MULTS_7_1(9)<=signed(MULTS_6_1(9)(PERCISION) & MULTS_6_1(9)(PERCISION downto 1))+signed(MULTS_6_2(9)(PERCISION) & MULTS_6_2(9)(PERCISION downto 1));



                        Enable_BIAS<='1';
		end if;


		------------------------------------STAGE-BIAS--------------------------------------
		if Enable_BIAS = '1' then

			BIAS_1<=(1+signed( MULTS_7_1(0)(PERCISION downto 1)));
			BIAS_2<=(1+signed( MULTS_7_1(1)(PERCISION downto 1)));
			BIAS_3<=(1+signed( MULTS_7_1(2)(PERCISION downto 1)));
			BIAS_4<=(1+signed( MULTS_7_1(3)(PERCISION downto 1)));
			BIAS_5<=(1+signed( MULTS_7_1(4)(PERCISION downto 1)));
			BIAS_6<=(1+signed( MULTS_7_1(5)(PERCISION downto 1)));
			BIAS_7<=(1+signed( MULTS_7_1(6)(PERCISION downto 1)));
			BIAS_8<=(1+signed( MULTS_7_1(7)(PERCISION downto 1)));
			BIAS_9<=(1+signed( MULTS_7_1(8)(PERCISION downto 1)));
			BIAS_10<=(1+signed( MULTS_7_1(9)(PERCISION downto 1)));

			Enable_ReLU<='1';
			
		end if;

		if SIG_STRIDE>1 and Enable_ReLU='1' then
                 SIG_STRIDE<=SIG_STRIDE-1; end if;

	if  Enable_ReLU='1' then
		if VALID_NXTLYR_PIX<VALID_LOCAL_PIX and SIG_STRIDE>(STRIDE-1) then

			if BIAS_1>0 then
			ReLU_1<=BIAS_1;
			DOUT_BUF_1_8<=std_logic_vector(BIAS_1);
			else
			ReLU_1<= (others => '0');
			DOUT_BUF_1_8<=(others => '0');
			end if;
			if BIAS_2>0 then
			ReLU_2<=BIAS_2;
			DOUT_BUF_2_8<=std_logic_vector(BIAS_2);
			else
			ReLU_2<= (others => '0');
			DOUT_BUF_2_8<=(others => '0');
			end if;
			if BIAS_3>0 then
			ReLU_3<=BIAS_3;
			DOUT_BUF_3_8<=std_logic_vector(BIAS_3);
			else
			ReLU_3<= (others => '0');
			DOUT_BUF_3_8<=(others => '0');
			end if;
			if BIAS_4>0 then
			ReLU_4<=BIAS_4;
			DOUT_BUF_4_8<=std_logic_vector(BIAS_4);
			else
			ReLU_4<= (others => '0');
			DOUT_BUF_4_8<=(others => '0');
			end if;
			if BIAS_5>0 then
			ReLU_5<=BIAS_5;
			DOUT_BUF_5_8<=std_logic_vector(BIAS_5);
			else
			ReLU_5<= (others => '0');
			DOUT_BUF_5_8<=(others => '0');
			end if;
			if BIAS_6>0 then
			ReLU_6<=BIAS_6;
			DOUT_BUF_6_8<=std_logic_vector(BIAS_6);
			else
			ReLU_6<= (others => '0');
			DOUT_BUF_6_8<=(others => '0');
			end if;
			if BIAS_7>0 then
			ReLU_7<=BIAS_7;
			DOUT_BUF_7_8<=std_logic_vector(BIAS_7);
			else
			ReLU_7<= (others => '0');
			DOUT_BUF_7_8<=(others => '0');
			end if;
			if BIAS_8>0 then
			ReLU_8<=BIAS_8;
			DOUT_BUF_8_8<=std_logic_vector(BIAS_8);
			else
			ReLU_8<= (others => '0');
			DOUT_BUF_8_8<=(others => '0');
			end if;
			if BIAS_9>0 then
			ReLU_9<=BIAS_9;
			DOUT_BUF_9_8<=std_logic_vector(BIAS_9);
			else
			ReLU_9<= (others => '0');
			DOUT_BUF_9_8<=(others => '0');
			end if;
			if BIAS_10>0 then
			ReLU_10<=BIAS_10;
			DOUT_BUF_10_8<=std_logic_vector(BIAS_10);
			else
			ReLU_10<= (others => '0');
			DOUT_BUF_10_8<=(others => '0');
			end if;

			EN_NXT_LYR_8<='1';FRST_TIM_EN_8<='1';
			OUT_PIXEL_COUNT<=OUT_PIXEL_COUNT+1;
		else
                       EN_NXT_LYR_8<='0';
                       DOUT_BUF_1_8<=(others => '0');
                       DOUT_BUF_2_8<=(others => '0');
                       DOUT_BUF_3_8<=(others => '0');
                       DOUT_BUF_4_8<=(others => '0');
                       DOUT_BUF_5_8<=(others => '0');
                       DOUT_BUF_6_8<=(others => '0');
                       DOUT_BUF_7_8<=(others => '0');
                       DOUT_BUF_8_8<=(others => '0');
                       DOUT_BUF_9_8<=(others => '0');
                       DOUT_BUF_10_8<=(others => '0');

		end if; -- VALIDPIXELS

		if VALID_NXTLYR_PIX=((VALID_LOCAL_PIX*STRIDE)-1) then VALID_NXTLYR_PIX<=0;SIG_STRIDE<=STRIDE;   -- reset sride and valid pixels
		else VALID_NXTLYR_PIX<=VALID_NXTLYR_PIX+1;end if; 

	end if;  --ReLU
elsif OUT_PIXEL_COUNT>=VALID_CYCLES  then INTERNAL_RST<='1';SIG_STRIDE<=STRIDE;EN_NXT_LYR_8<='1';  -- order is very important
else  EN_NXT_LYR_8<='0';-- In case stream stopped

end if; -- end enable 
end if; -- for RST	
end if; -- rising edge
end process LAYER_8;

DOUT_1_8<=DOUT_BUF_1_8;
DOUT_2_8<=DOUT_BUF_2_8;
DOUT_3_8<=DOUT_BUF_3_8;
DOUT_4_8<=DOUT_BUF_4_8;
DOUT_5_8<=DOUT_BUF_5_8;
DOUT_6_8<=DOUT_BUF_6_8;
DOUT_7_8<=DOUT_BUF_7_8;
DOUT_8_8<=DOUT_BUF_8_8;
DOUT_9_8<=DOUT_BUF_9_8;
DOUT_10_8<=DOUT_BUF_10_8;

end Behavioral;
------------------------------ ARCHITECTURE DECLARATION - END---------------------------------------------

