------------------------------------------HEADER START"------------------------------------------
--THIS FILE WAS GENERATED USING HIGH LANGUAGE DESCRIPTION TOOL DESIGNED BY: MUHAMMAD HAMDAN
--TOOL VERSION: 0.1
--GENERATION DATE/TIME:Mon Apr 06 09:42:53 CDT 2020
------------------------------------------HEADER END"--------------------------------------------



------------------------------DESCRIPTION AND LIBRARY DECLARATION-START---------------------------
-- Engineer:       Muhammad Hamdan
-- Design Name:    HDL GENERATION - CONV LAYER 
-- Module Name:    FC - Behavioral 
-- Project Name:   CNN accelerator
-- Number of Total Operaiton: 336
-- Number of Clock Cycles: 48
-- Number of GOPS = 3.0
-------------------------------------------------Total Number of Operations for the Entire Model:10
-- Target Devices: Zynq-XC7Z020
-- Description: 
-- Dependencies: 
-- Revision:0.010 


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_arith.all;

entity FC_LAYER_7 is

GENERIC
 	( 
	constant PERCISION      : positive := 5; 	
	constant DOUT_WIDTH     : positive := 5; 	
	constant BIAS_SIZE      : positive := 5;
	constant MULT_SIZE      : positive := 10;
	constant BASE_DIN_WIDTH : positive := 62;
	constant DIN_WIDTH      : positive := 5;
	constant IMAGE_WIDTH    : positive := 1;
	constant IMAGE_SIZE     : positive := 1024;	
	constant F_SIZE         : positive := 1;
	constant PF_X2_SIZE     : positive := 25;
	constant WEIGHT_SIZE    : positive := 5;
	constant BIASES_SIZE	: positive := 2;
	constant PADDING        : positive := 1;
	constant STRIDE         : positive := 1;
	constant FEATURE_MAPS   : positive := 84;
	constant VALID_CYCLES   : positive := 25;
	constant VALID_LOCAL_PIX: positive := 5;
	constant ADD_TREE_DEPTH : positive := 1;
	constant INPUT_DEPTH    : positive := 7;
	constant INNER_PXL_SUM  : positive := 1;
	constant SUM_PEXILS     : positive := 87;
	constant MULT_SUM_D_1   : positive := 60;
	constant MULT_SUM_SIZE_1: positive := 6;
	constant MULT_SUM_D_2   : positive := 30;
	constant MULT_SUM_SIZE_2: positive := 6;
	constant MULT_SUM_D_3   : positive := 15;
	constant MULT_SUM_SIZE_3: positive := 6;
	constant MULT_SUM_D_4   : positive := 8;
	constant MULT_SUM_SIZE_4: positive := 6;
	constant MULT_SUM_D_5   : positive := 4;
	constant MULT_SUM_SIZE_5: positive := 6;
	constant MULT_SUM_D_6   : positive := 2;
	constant MULT_SUM_SIZE_6: positive := 6;
	constant MULT_SUM_D_7   : positive := 1;
	constant MULT_SUM_SIZE_7: positive := 6;
	constant LOCAL_OUTPUT   : positive := 5	
		); 

port(
	DIN_1_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_2_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_3_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_4_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_5_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_6_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_7_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_8_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_9_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_10_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_11_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_12_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_13_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_14_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_15_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_16_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_17_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_18_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_19_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_20_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_21_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_22_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_23_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_24_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_25_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_26_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_27_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_28_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_29_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_30_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_31_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_32_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_33_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_34_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_35_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_36_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_37_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_38_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_39_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_40_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_41_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_42_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_43_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_44_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_45_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_46_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_47_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_48_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_49_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_50_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_51_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_52_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_53_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_54_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_55_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_56_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_57_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_58_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_59_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_60_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_61_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_62_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_63_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_64_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_65_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_66_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_67_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_68_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_69_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_70_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_71_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_72_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_73_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_74_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_75_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_76_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_77_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_78_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_79_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_80_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_81_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_82_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_83_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_84_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_85_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_86_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_87_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_88_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_89_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_90_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_91_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_92_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_93_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_94_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_95_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_96_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_97_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_98_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_99_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_100_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_101_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_102_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_103_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_104_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_105_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_106_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_107_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_108_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_109_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_110_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_111_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_112_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_113_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_114_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_115_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_116_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_117_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_118_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_119_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_120_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	CLK,RST         :IN std_logic;
   	DIS_STREAM      :OUT std_logic; 				-- S_AXIS_TVALID  : Data in is valid
   	EN_STREAM       :IN std_logic; 					-- S_AXIS_TREADY  : Ready to accept data in 
	EN_STREAM_OUT_7 :OUT std_logic; 			-- M_AXIS_TREADY  : Connected slave device is ready to accept data out/ Internal Enable
	VALID_OUT_7     :OUT std_logic;                         -- M_AXIS_TVALID  : Data out is valid
	EN_LOC_STREAM_7 :IN std_logic;
	DOUT_1_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_2_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_3_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_4_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_5_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_6_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_7_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_8_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_9_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_10_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	INTERNAL_RST    :OUT std_logic
	);	

end FC_LAYER_7;

------------------------------ ARCHITECTURE DECLARATION - START---------------------------------------------

architecture Behavioral of FC_LAYER_7 is

------------------------------ INTERNAL FIXED CONSTANT & SIGNALS DECLARATION - START---------------------------------------------
type       FILTER_TYPE             is array (0 to PF_X2_SIZE-1) of signed(WEIGHT_SIZE- 1 downto 0);
signal     VALID_NXTLYR_PIX        :integer range 0 to VALID_CYCLES;
signal     PIXEL_COUNT             :integer range 0 to VALID_CYCLES;
signal     OUT_PIXEL_COUNT         :integer range 0 to VALID_CYCLES;
signal     EN_NXT_LYR_7            :std_logic;
signal     FRST_TIM_EN_7           :std_logic;
signal     Enable_MULT             :std_logic;
signal     Enable_ADDER            :std_logic;
signal     Enable_ReLU             :std_logic;
signal     Enable_BIAS             :std_logic;
signal     COUNT_PIX               :integer range 0 to PF_X2_SIZE;
signal     SIG_STRIDE              :integer range 0 to IMAGE_SIZE;
signal     PADDING_count           :integer range 0 to IMAGE_SIZE; -- TEMPORARY
signal     ROW_COUNT               :integer range 0 to IMAGE_SIZE; -- TEMPORARY


------------------------------ INTERNAL DYNAMIC SIGNALS DECLARATION ARRAY TYPE- START---------------------------------------------


type   MULT_X		is array (0 to FEATURE_MAPS-1) of signed(MULT_SIZE- 1 downto 0);
signal MULT_1:MULT_X;
signal MULT_2:MULT_X;
signal MULT_3:MULT_X;
signal MULT_4:MULT_X;
signal MULT_5:MULT_X;
signal MULT_6:MULT_X;
signal MULT_7:MULT_X;
signal MULT_8:MULT_X;
signal MULT_9:MULT_X;
signal MULT_10:MULT_X;
signal MULT_11:MULT_X;
signal MULT_12:MULT_X;
signal MULT_13:MULT_X;
signal MULT_14:MULT_X;
signal MULT_15:MULT_X;
signal MULT_16:MULT_X;
signal MULT_17:MULT_X;
signal MULT_18:MULT_X;
signal MULT_19:MULT_X;
signal MULT_20:MULT_X;
signal MULT_21:MULT_X;
signal MULT_22:MULT_X;
signal MULT_23:MULT_X;
signal MULT_24:MULT_X;
signal MULT_25:MULT_X;
signal MULT_26:MULT_X;
signal MULT_27:MULT_X;
signal MULT_28:MULT_X;
signal MULT_29:MULT_X;
signal MULT_30:MULT_X;
signal MULT_31:MULT_X;
signal MULT_32:MULT_X;
signal MULT_33:MULT_X;
signal MULT_34:MULT_X;
signal MULT_35:MULT_X;
signal MULT_36:MULT_X;
signal MULT_37:MULT_X;
signal MULT_38:MULT_X;
signal MULT_39:MULT_X;
signal MULT_40:MULT_X;
signal MULT_41:MULT_X;
signal MULT_42:MULT_X;
signal MULT_43:MULT_X;
signal MULT_44:MULT_X;
signal MULT_45:MULT_X;
signal MULT_46:MULT_X;
signal MULT_47:MULT_X;
signal MULT_48:MULT_X;
signal MULT_49:MULT_X;
signal MULT_50:MULT_X;
signal MULT_51:MULT_X;
signal MULT_52:MULT_X;
signal MULT_53:MULT_X;
signal MULT_54:MULT_X;
signal MULT_55:MULT_X;
signal MULT_56:MULT_X;
signal MULT_57:MULT_X;
signal MULT_58:MULT_X;
signal MULT_59:MULT_X;
signal MULT_60:MULT_X;
signal MULT_61:MULT_X;
signal MULT_62:MULT_X;
signal MULT_63:MULT_X;
signal MULT_64:MULT_X;
signal MULT_65:MULT_X;
signal MULT_66:MULT_X;
signal MULT_67:MULT_X;
signal MULT_68:MULT_X;
signal MULT_69:MULT_X;
signal MULT_70:MULT_X;
signal MULT_71:MULT_X;
signal MULT_72:MULT_X;
signal MULT_73:MULT_X;
signal MULT_74:MULT_X;
signal MULT_75:MULT_X;
signal MULT_76:MULT_X;
signal MULT_77:MULT_X;
signal MULT_78:MULT_X;
signal MULT_79:MULT_X;
signal MULT_80:MULT_X;
signal MULT_81:MULT_X;
signal MULT_82:MULT_X;
signal MULT_83:MULT_X;
signal MULT_84:MULT_X;
signal MULT_85:MULT_X;
signal MULT_86:MULT_X;
signal MULT_87:MULT_X;
signal MULT_88:MULT_X;
signal MULT_89:MULT_X;
signal MULT_90:MULT_X;
signal MULT_91:MULT_X;
signal MULT_92:MULT_X;
signal MULT_93:MULT_X;
signal MULT_94:MULT_X;
signal MULT_95:MULT_X;
signal MULT_96:MULT_X;
signal MULT_97:MULT_X;
signal MULT_98:MULT_X;
signal MULT_99:MULT_X;
signal MULT_100:MULT_X;
signal MULT_101:MULT_X;
signal MULT_102:MULT_X;
signal MULT_103:MULT_X;
signal MULT_104:MULT_X;
signal MULT_105:MULT_X;
signal MULT_106:MULT_X;
signal MULT_107:MULT_X;
signal MULT_108:MULT_X;
signal MULT_109:MULT_X;
signal MULT_110:MULT_X;
signal MULT_111:MULT_X;
signal MULT_112:MULT_X;
signal MULT_113:MULT_X;
signal MULT_114:MULT_X;
signal MULT_115:MULT_X;
signal MULT_116:MULT_X;
signal MULT_117:MULT_X;
signal MULT_118:MULT_X;
signal MULT_119:MULT_X;
signal MULT_120:MULT_X;
signal DOUT_BUF_1_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_1		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_1		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_2_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_2		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_2		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_3_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_3		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_3		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_4_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_4		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_4		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_5_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_5		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_5		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_6_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_6		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_6		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_7_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_7		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_7		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_8_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_8		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_8		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_9_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_9		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_9		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_10_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_10		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_10		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_11_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_11		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_11		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_12_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_12		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_12		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_13_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_13		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_13		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_14_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_14		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_14		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_15_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_15		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_15		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_16_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_16		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_16		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_17_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_17		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_17		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_18_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_18		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_18		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_19_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_19		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_19		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_20_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_20		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_20		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_21_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_21		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_21		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_22_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_22		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_22		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_23_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_23		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_23		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_24_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_24		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_24		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_25_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_25		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_25		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_26_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_26		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_26		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_27_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_27		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_27		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_28_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_28		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_28		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_29_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_29		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_29		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_30_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_30		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_30		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_31_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_31		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_31		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_32_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_32		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_32		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_33_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_33		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_33		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_34_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_34		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_34		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_35_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_35		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_35		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_36_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_36		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_36		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_37_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_37		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_37		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_38_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_38		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_38		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_39_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_39		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_39		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_40_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_40		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_40		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_41_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_41		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_41		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_42_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_42		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_42		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_43_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_43		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_43		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_44_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_44		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_44		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_45_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_45		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_45		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_46_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_46		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_46		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_47_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_47		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_47		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_48_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_48		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_48		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_49_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_49		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_49		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_50_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_50		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_50		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_51_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_51		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_51		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_52_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_52		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_52		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_53_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_53		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_53		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_54_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_54		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_54		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_55_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_55		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_55		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_56_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_56		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_56		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_57_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_57		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_57		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_58_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_58		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_58		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_59_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_59		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_59		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_60_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_60		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_60		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_61_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_61		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_61		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_62_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_62		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_62		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_63_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_63		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_63		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_64_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_64		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_64		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_65_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_65		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_65		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_66_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_66		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_66		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_67_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_67		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_67		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_68_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_68		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_68		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_69_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_69		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_69		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_70_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_70		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_70		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_71_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_71		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_71		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_72_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_72		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_72		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_73_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_73		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_73		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_74_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_74		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_74		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_75_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_75		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_75		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_76_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_76		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_76		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_77_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_77		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_77		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_78_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_78		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_78		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_79_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_79		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_79		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_80_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_80		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_80		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_81_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_81		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_81		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_82_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_82		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_82		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_83_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_83		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_83		: signed(BIAS_SIZE-1   downto 0);
signal DOUT_BUF_84_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_84		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_84		: signed(BIAS_SIZE-1   downto 0);


------------------------------------------------------ MULT SUMMATION DECLARATION-----------------------------------------------------------
signal SUM_PIXELS_1: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_2: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_3: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_4: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_5: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_6: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_7: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_8: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_9: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_10: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_11: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_12: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_13: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_14: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_15: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_16: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_17: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_18: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_19: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_20: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_21: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_22: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_23: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_24: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_25: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_26: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_27: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_28: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_29: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_30: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_31: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_32: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_33: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_34: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_35: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_36: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_37: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_38: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_39: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_40: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_41: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_42: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_43: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_44: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_45: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_46: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_47: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_48: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_49: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_50: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_51: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_52: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_53: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_54: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_55: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_56: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_57: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_58: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_59: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_60: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_61: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_62: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_63: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_64: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_65: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_66: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_67: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_68: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_69: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_70: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_71: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_72: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_73: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_74: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_75: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_76: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_77: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_78: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_79: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_80: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_81: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_82: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_83: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_84: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_85: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_86: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_87: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_88: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_89: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_90: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_91: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_92: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_93: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_94: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_95: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_96: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_97: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_98: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_99: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_100: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_101: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_102: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_103: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_104: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_105: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_106: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_107: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_108: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_109: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_110: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_111: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_112: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_113: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_114: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_115: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_116: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_117: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_118: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_119: signed(SUM_PEXILS-1 downto 0);
signal SUM_PIXELS_120: signed(SUM_PEXILS-1 downto 0);
type    MULT_X_SUM_1	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_1- 1 downto 0);
signal  EN_SUM_MULT_1	: std_logic;
signal  MULTS_1_1:MULT_X_SUM_1;
signal  MULTS_1_2:MULT_X_SUM_1;
signal  MULTS_1_3:MULT_X_SUM_1;
signal  MULTS_1_4:MULT_X_SUM_1;
signal  MULTS_1_5:MULT_X_SUM_1;
signal  MULTS_1_6:MULT_X_SUM_1;
signal  MULTS_1_7:MULT_X_SUM_1;
signal  MULTS_1_8:MULT_X_SUM_1;
signal  MULTS_1_9:MULT_X_SUM_1;
signal  MULTS_1_10:MULT_X_SUM_1;
signal  MULTS_1_11:MULT_X_SUM_1;
signal  MULTS_1_12:MULT_X_SUM_1;
signal  MULTS_1_13:MULT_X_SUM_1;
signal  MULTS_1_14:MULT_X_SUM_1;
signal  MULTS_1_15:MULT_X_SUM_1;
signal  MULTS_1_16:MULT_X_SUM_1;
signal  MULTS_1_17:MULT_X_SUM_1;
signal  MULTS_1_18:MULT_X_SUM_1;
signal  MULTS_1_19:MULT_X_SUM_1;
signal  MULTS_1_20:MULT_X_SUM_1;
signal  MULTS_1_21:MULT_X_SUM_1;
signal  MULTS_1_22:MULT_X_SUM_1;
signal  MULTS_1_23:MULT_X_SUM_1;
signal  MULTS_1_24:MULT_X_SUM_1;
signal  MULTS_1_25:MULT_X_SUM_1;
signal  MULTS_1_26:MULT_X_SUM_1;
signal  MULTS_1_27:MULT_X_SUM_1;
signal  MULTS_1_28:MULT_X_SUM_1;
signal  MULTS_1_29:MULT_X_SUM_1;
signal  MULTS_1_30:MULT_X_SUM_1;
signal  MULTS_1_31:MULT_X_SUM_1;
signal  MULTS_1_32:MULT_X_SUM_1;
signal  MULTS_1_33:MULT_X_SUM_1;
signal  MULTS_1_34:MULT_X_SUM_1;
signal  MULTS_1_35:MULT_X_SUM_1;
signal  MULTS_1_36:MULT_X_SUM_1;
signal  MULTS_1_37:MULT_X_SUM_1;
signal  MULTS_1_38:MULT_X_SUM_1;
signal  MULTS_1_39:MULT_X_SUM_1;
signal  MULTS_1_40:MULT_X_SUM_1;
signal  MULTS_1_41:MULT_X_SUM_1;
signal  MULTS_1_42:MULT_X_SUM_1;
signal  MULTS_1_43:MULT_X_SUM_1;
signal  MULTS_1_44:MULT_X_SUM_1;
signal  MULTS_1_45:MULT_X_SUM_1;
signal  MULTS_1_46:MULT_X_SUM_1;
signal  MULTS_1_47:MULT_X_SUM_1;
signal  MULTS_1_48:MULT_X_SUM_1;
signal  MULTS_1_49:MULT_X_SUM_1;
signal  MULTS_1_50:MULT_X_SUM_1;
signal  MULTS_1_51:MULT_X_SUM_1;
signal  MULTS_1_52:MULT_X_SUM_1;
signal  MULTS_1_53:MULT_X_SUM_1;
signal  MULTS_1_54:MULT_X_SUM_1;
signal  MULTS_1_55:MULT_X_SUM_1;
signal  MULTS_1_56:MULT_X_SUM_1;
signal  MULTS_1_57:MULT_X_SUM_1;
signal  MULTS_1_58:MULT_X_SUM_1;
signal  MULTS_1_59:MULT_X_SUM_1;
signal  MULTS_1_60:MULT_X_SUM_1;
signal  MULTS_1_61:MULT_X_SUM_1;
signal  MULTS_1_62:MULT_X_SUM_1;
signal  MULTS_1_63:MULT_X_SUM_1;
signal  MULTS_1_64:MULT_X_SUM_1;
signal  MULTS_1_65:MULT_X_SUM_1;
signal  MULTS_1_66:MULT_X_SUM_1;
signal  MULTS_1_67:MULT_X_SUM_1;
signal  MULTS_1_68:MULT_X_SUM_1;
signal  MULTS_1_69:MULT_X_SUM_1;
signal  MULTS_1_70:MULT_X_SUM_1;
signal  MULTS_1_71:MULT_X_SUM_1;
signal  MULTS_1_72:MULT_X_SUM_1;
signal  MULTS_1_73:MULT_X_SUM_1;
signal  MULTS_1_74:MULT_X_SUM_1;
signal  MULTS_1_75:MULT_X_SUM_1;
signal  MULTS_1_76:MULT_X_SUM_1;
signal  MULTS_1_77:MULT_X_SUM_1;
signal  MULTS_1_78:MULT_X_SUM_1;
signal  MULTS_1_79:MULT_X_SUM_1;
signal  MULTS_1_80:MULT_X_SUM_1;
signal  MULTS_1_81:MULT_X_SUM_1;
signal  MULTS_1_82:MULT_X_SUM_1;
signal  MULTS_1_83:MULT_X_SUM_1;
signal  MULTS_1_84:MULT_X_SUM_1;
signal  MULTS_1_85:MULT_X_SUM_1;
signal  MULTS_1_86:MULT_X_SUM_1;
signal  MULTS_1_87:MULT_X_SUM_1;
signal  MULTS_1_88:MULT_X_SUM_1;
signal  MULTS_1_89:MULT_X_SUM_1;
signal  MULTS_1_90:MULT_X_SUM_1;
signal  MULTS_1_91:MULT_X_SUM_1;
signal  MULTS_1_92:MULT_X_SUM_1;
signal  MULTS_1_93:MULT_X_SUM_1;
signal  MULTS_1_94:MULT_X_SUM_1;
signal  MULTS_1_95:MULT_X_SUM_1;
signal  MULTS_1_96:MULT_X_SUM_1;
signal  MULTS_1_97:MULT_X_SUM_1;
signal  MULTS_1_98:MULT_X_SUM_1;
signal  MULTS_1_99:MULT_X_SUM_1;
signal  MULTS_1_100:MULT_X_SUM_1;
signal  MULTS_1_101:MULT_X_SUM_1;
signal  MULTS_1_102:MULT_X_SUM_1;
signal  MULTS_1_103:MULT_X_SUM_1;
signal  MULTS_1_104:MULT_X_SUM_1;
signal  MULTS_1_105:MULT_X_SUM_1;
signal  MULTS_1_106:MULT_X_SUM_1;
signal  MULTS_1_107:MULT_X_SUM_1;
signal  MULTS_1_108:MULT_X_SUM_1;
signal  MULTS_1_109:MULT_X_SUM_1;
signal  MULTS_1_110:MULT_X_SUM_1;
signal  MULTS_1_111:MULT_X_SUM_1;
signal  MULTS_1_112:MULT_X_SUM_1;
signal  MULTS_1_113:MULT_X_SUM_1;
signal  MULTS_1_114:MULT_X_SUM_1;
signal  MULTS_1_115:MULT_X_SUM_1;
signal  MULTS_1_116:MULT_X_SUM_1;
signal  MULTS_1_117:MULT_X_SUM_1;
signal  MULTS_1_118:MULT_X_SUM_1;
signal  MULTS_1_119:MULT_X_SUM_1;
signal  MULTS_1_120:MULT_X_SUM_1;
type    MULT_X_SUM_2	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_2- 1 downto 0);
signal  EN_SUM_MULT_2	: std_logic;
signal  MULTS_2_1:MULT_X_SUM_2;
signal  MULTS_2_2:MULT_X_SUM_2;
signal  MULTS_2_3:MULT_X_SUM_2;
signal  MULTS_2_4:MULT_X_SUM_2;
signal  MULTS_2_5:MULT_X_SUM_2;
signal  MULTS_2_6:MULT_X_SUM_2;
signal  MULTS_2_7:MULT_X_SUM_2;
signal  MULTS_2_8:MULT_X_SUM_2;
signal  MULTS_2_9:MULT_X_SUM_2;
signal  MULTS_2_10:MULT_X_SUM_2;
signal  MULTS_2_11:MULT_X_SUM_2;
signal  MULTS_2_12:MULT_X_SUM_2;
signal  MULTS_2_13:MULT_X_SUM_2;
signal  MULTS_2_14:MULT_X_SUM_2;
signal  MULTS_2_15:MULT_X_SUM_2;
signal  MULTS_2_16:MULT_X_SUM_2;
signal  MULTS_2_17:MULT_X_SUM_2;
signal  MULTS_2_18:MULT_X_SUM_2;
signal  MULTS_2_19:MULT_X_SUM_2;
signal  MULTS_2_20:MULT_X_SUM_2;
signal  MULTS_2_21:MULT_X_SUM_2;
signal  MULTS_2_22:MULT_X_SUM_2;
signal  MULTS_2_23:MULT_X_SUM_2;
signal  MULTS_2_24:MULT_X_SUM_2;
signal  MULTS_2_25:MULT_X_SUM_2;
signal  MULTS_2_26:MULT_X_SUM_2;
signal  MULTS_2_27:MULT_X_SUM_2;
signal  MULTS_2_28:MULT_X_SUM_2;
signal  MULTS_2_29:MULT_X_SUM_2;
signal  MULTS_2_30:MULT_X_SUM_2;
signal  MULTS_2_31:MULT_X_SUM_2;
signal  MULTS_2_32:MULT_X_SUM_2;
signal  MULTS_2_33:MULT_X_SUM_2;
signal  MULTS_2_34:MULT_X_SUM_2;
signal  MULTS_2_35:MULT_X_SUM_2;
signal  MULTS_2_36:MULT_X_SUM_2;
signal  MULTS_2_37:MULT_X_SUM_2;
signal  MULTS_2_38:MULT_X_SUM_2;
signal  MULTS_2_39:MULT_X_SUM_2;
signal  MULTS_2_40:MULT_X_SUM_2;
signal  MULTS_2_41:MULT_X_SUM_2;
signal  MULTS_2_42:MULT_X_SUM_2;
signal  MULTS_2_43:MULT_X_SUM_2;
signal  MULTS_2_44:MULT_X_SUM_2;
signal  MULTS_2_45:MULT_X_SUM_2;
signal  MULTS_2_46:MULT_X_SUM_2;
signal  MULTS_2_47:MULT_X_SUM_2;
signal  MULTS_2_48:MULT_X_SUM_2;
signal  MULTS_2_49:MULT_X_SUM_2;
signal  MULTS_2_50:MULT_X_SUM_2;
signal  MULTS_2_51:MULT_X_SUM_2;
signal  MULTS_2_52:MULT_X_SUM_2;
signal  MULTS_2_53:MULT_X_SUM_2;
signal  MULTS_2_54:MULT_X_SUM_2;
signal  MULTS_2_55:MULT_X_SUM_2;
signal  MULTS_2_56:MULT_X_SUM_2;
signal  MULTS_2_57:MULT_X_SUM_2;
signal  MULTS_2_58:MULT_X_SUM_2;
signal  MULTS_2_59:MULT_X_SUM_2;
signal  MULTS_2_60:MULT_X_SUM_2;
signal  MULTS_2_61:MULT_X_SUM_2;
signal  MULTS_2_62:MULT_X_SUM_2;
signal  MULTS_2_63:MULT_X_SUM_2;
signal  MULTS_2_64:MULT_X_SUM_2;
signal  MULTS_2_65:MULT_X_SUM_2;
signal  MULTS_2_66:MULT_X_SUM_2;
signal  MULTS_2_67:MULT_X_SUM_2;
signal  MULTS_2_68:MULT_X_SUM_2;
signal  MULTS_2_69:MULT_X_SUM_2;
signal  MULTS_2_70:MULT_X_SUM_2;
signal  MULTS_2_71:MULT_X_SUM_2;
signal  MULTS_2_72:MULT_X_SUM_2;
signal  MULTS_2_73:MULT_X_SUM_2;
signal  MULTS_2_74:MULT_X_SUM_2;
signal  MULTS_2_75:MULT_X_SUM_2;
signal  MULTS_2_76:MULT_X_SUM_2;
signal  MULTS_2_77:MULT_X_SUM_2;
signal  MULTS_2_78:MULT_X_SUM_2;
signal  MULTS_2_79:MULT_X_SUM_2;
signal  MULTS_2_80:MULT_X_SUM_2;
signal  MULTS_2_81:MULT_X_SUM_2;
signal  MULTS_2_82:MULT_X_SUM_2;
signal  MULTS_2_83:MULT_X_SUM_2;
signal  MULTS_2_84:MULT_X_SUM_2;
signal  MULTS_2_85:MULT_X_SUM_2;
signal  MULTS_2_86:MULT_X_SUM_2;
signal  MULTS_2_87:MULT_X_SUM_2;
signal  MULTS_2_88:MULT_X_SUM_2;
signal  MULTS_2_89:MULT_X_SUM_2;
signal  MULTS_2_90:MULT_X_SUM_2;
signal  MULTS_2_91:MULT_X_SUM_2;
signal  MULTS_2_92:MULT_X_SUM_2;
signal  MULTS_2_93:MULT_X_SUM_2;
signal  MULTS_2_94:MULT_X_SUM_2;
signal  MULTS_2_95:MULT_X_SUM_2;
signal  MULTS_2_96:MULT_X_SUM_2;
signal  MULTS_2_97:MULT_X_SUM_2;
signal  MULTS_2_98:MULT_X_SUM_2;
signal  MULTS_2_99:MULT_X_SUM_2;
signal  MULTS_2_100:MULT_X_SUM_2;
signal  MULTS_2_101:MULT_X_SUM_2;
signal  MULTS_2_102:MULT_X_SUM_2;
signal  MULTS_2_103:MULT_X_SUM_2;
signal  MULTS_2_104:MULT_X_SUM_2;
signal  MULTS_2_105:MULT_X_SUM_2;
signal  MULTS_2_106:MULT_X_SUM_2;
signal  MULTS_2_107:MULT_X_SUM_2;
signal  MULTS_2_108:MULT_X_SUM_2;
signal  MULTS_2_109:MULT_X_SUM_2;
signal  MULTS_2_110:MULT_X_SUM_2;
signal  MULTS_2_111:MULT_X_SUM_2;
signal  MULTS_2_112:MULT_X_SUM_2;
signal  MULTS_2_113:MULT_X_SUM_2;
signal  MULTS_2_114:MULT_X_SUM_2;
signal  MULTS_2_115:MULT_X_SUM_2;
signal  MULTS_2_116:MULT_X_SUM_2;
signal  MULTS_2_117:MULT_X_SUM_2;
signal  MULTS_2_118:MULT_X_SUM_2;
signal  MULTS_2_119:MULT_X_SUM_2;
signal  MULTS_2_120:MULT_X_SUM_2;
type    MULT_X_SUM_3	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_3- 1 downto 0);
signal  EN_SUM_MULT_3	: std_logic;
signal  MULTS_3_1:MULT_X_SUM_3;
signal  MULTS_3_2:MULT_X_SUM_3;
signal  MULTS_3_3:MULT_X_SUM_3;
signal  MULTS_3_4:MULT_X_SUM_3;
signal  MULTS_3_5:MULT_X_SUM_3;
signal  MULTS_3_6:MULT_X_SUM_3;
signal  MULTS_3_7:MULT_X_SUM_3;
signal  MULTS_3_8:MULT_X_SUM_3;
signal  MULTS_3_9:MULT_X_SUM_3;
signal  MULTS_3_10:MULT_X_SUM_3;
signal  MULTS_3_11:MULT_X_SUM_3;
signal  MULTS_3_12:MULT_X_SUM_3;
signal  MULTS_3_13:MULT_X_SUM_3;
signal  MULTS_3_14:MULT_X_SUM_3;
signal  MULTS_3_15:MULT_X_SUM_3;
signal  MULTS_3_16:MULT_X_SUM_3;
signal  MULTS_3_17:MULT_X_SUM_3;
signal  MULTS_3_18:MULT_X_SUM_3;
signal  MULTS_3_19:MULT_X_SUM_3;
signal  MULTS_3_20:MULT_X_SUM_3;
signal  MULTS_3_21:MULT_X_SUM_3;
signal  MULTS_3_22:MULT_X_SUM_3;
signal  MULTS_3_23:MULT_X_SUM_3;
signal  MULTS_3_24:MULT_X_SUM_3;
signal  MULTS_3_25:MULT_X_SUM_3;
signal  MULTS_3_26:MULT_X_SUM_3;
signal  MULTS_3_27:MULT_X_SUM_3;
signal  MULTS_3_28:MULT_X_SUM_3;
signal  MULTS_3_29:MULT_X_SUM_3;
signal  MULTS_3_30:MULT_X_SUM_3;
signal  MULTS_3_31:MULT_X_SUM_3;
signal  MULTS_3_32:MULT_X_SUM_3;
signal  MULTS_3_33:MULT_X_SUM_3;
signal  MULTS_3_34:MULT_X_SUM_3;
signal  MULTS_3_35:MULT_X_SUM_3;
signal  MULTS_3_36:MULT_X_SUM_3;
signal  MULTS_3_37:MULT_X_SUM_3;
signal  MULTS_3_38:MULT_X_SUM_3;
signal  MULTS_3_39:MULT_X_SUM_3;
signal  MULTS_3_40:MULT_X_SUM_3;
signal  MULTS_3_41:MULT_X_SUM_3;
signal  MULTS_3_42:MULT_X_SUM_3;
signal  MULTS_3_43:MULT_X_SUM_3;
signal  MULTS_3_44:MULT_X_SUM_3;
signal  MULTS_3_45:MULT_X_SUM_3;
signal  MULTS_3_46:MULT_X_SUM_3;
signal  MULTS_3_47:MULT_X_SUM_3;
signal  MULTS_3_48:MULT_X_SUM_3;
signal  MULTS_3_49:MULT_X_SUM_3;
signal  MULTS_3_50:MULT_X_SUM_3;
signal  MULTS_3_51:MULT_X_SUM_3;
signal  MULTS_3_52:MULT_X_SUM_3;
signal  MULTS_3_53:MULT_X_SUM_3;
signal  MULTS_3_54:MULT_X_SUM_3;
signal  MULTS_3_55:MULT_X_SUM_3;
signal  MULTS_3_56:MULT_X_SUM_3;
signal  MULTS_3_57:MULT_X_SUM_3;
signal  MULTS_3_58:MULT_X_SUM_3;
signal  MULTS_3_59:MULT_X_SUM_3;
signal  MULTS_3_60:MULT_X_SUM_3;
signal  MULTS_3_61:MULT_X_SUM_3;
signal  MULTS_3_62:MULT_X_SUM_3;
signal  MULTS_3_63:MULT_X_SUM_3;
signal  MULTS_3_64:MULT_X_SUM_3;
signal  MULTS_3_65:MULT_X_SUM_3;
signal  MULTS_3_66:MULT_X_SUM_3;
signal  MULTS_3_67:MULT_X_SUM_3;
signal  MULTS_3_68:MULT_X_SUM_3;
signal  MULTS_3_69:MULT_X_SUM_3;
signal  MULTS_3_70:MULT_X_SUM_3;
signal  MULTS_3_71:MULT_X_SUM_3;
signal  MULTS_3_72:MULT_X_SUM_3;
signal  MULTS_3_73:MULT_X_SUM_3;
signal  MULTS_3_74:MULT_X_SUM_3;
signal  MULTS_3_75:MULT_X_SUM_3;
signal  MULTS_3_76:MULT_X_SUM_3;
signal  MULTS_3_77:MULT_X_SUM_3;
signal  MULTS_3_78:MULT_X_SUM_3;
signal  MULTS_3_79:MULT_X_SUM_3;
signal  MULTS_3_80:MULT_X_SUM_3;
signal  MULTS_3_81:MULT_X_SUM_3;
signal  MULTS_3_82:MULT_X_SUM_3;
signal  MULTS_3_83:MULT_X_SUM_3;
signal  MULTS_3_84:MULT_X_SUM_3;
signal  MULTS_3_85:MULT_X_SUM_3;
signal  MULTS_3_86:MULT_X_SUM_3;
signal  MULTS_3_87:MULT_X_SUM_3;
signal  MULTS_3_88:MULT_X_SUM_3;
signal  MULTS_3_89:MULT_X_SUM_3;
signal  MULTS_3_90:MULT_X_SUM_3;
signal  MULTS_3_91:MULT_X_SUM_3;
signal  MULTS_3_92:MULT_X_SUM_3;
signal  MULTS_3_93:MULT_X_SUM_3;
signal  MULTS_3_94:MULT_X_SUM_3;
signal  MULTS_3_95:MULT_X_SUM_3;
signal  MULTS_3_96:MULT_X_SUM_3;
signal  MULTS_3_97:MULT_X_SUM_3;
signal  MULTS_3_98:MULT_X_SUM_3;
signal  MULTS_3_99:MULT_X_SUM_3;
signal  MULTS_3_100:MULT_X_SUM_3;
signal  MULTS_3_101:MULT_X_SUM_3;
signal  MULTS_3_102:MULT_X_SUM_3;
signal  MULTS_3_103:MULT_X_SUM_3;
signal  MULTS_3_104:MULT_X_SUM_3;
signal  MULTS_3_105:MULT_X_SUM_3;
signal  MULTS_3_106:MULT_X_SUM_3;
signal  MULTS_3_107:MULT_X_SUM_3;
signal  MULTS_3_108:MULT_X_SUM_3;
signal  MULTS_3_109:MULT_X_SUM_3;
signal  MULTS_3_110:MULT_X_SUM_3;
signal  MULTS_3_111:MULT_X_SUM_3;
signal  MULTS_3_112:MULT_X_SUM_3;
signal  MULTS_3_113:MULT_X_SUM_3;
signal  MULTS_3_114:MULT_X_SUM_3;
signal  MULTS_3_115:MULT_X_SUM_3;
signal  MULTS_3_116:MULT_X_SUM_3;
signal  MULTS_3_117:MULT_X_SUM_3;
signal  MULTS_3_118:MULT_X_SUM_3;
signal  MULTS_3_119:MULT_X_SUM_3;
signal  MULTS_3_120:MULT_X_SUM_3;
type    MULT_X_SUM_4	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_4- 1 downto 0);
signal  EN_SUM_MULT_4	: std_logic;
signal  MULTS_4_1:MULT_X_SUM_4;
signal  MULTS_4_2:MULT_X_SUM_4;
signal  MULTS_4_3:MULT_X_SUM_4;
signal  MULTS_4_4:MULT_X_SUM_4;
signal  MULTS_4_5:MULT_X_SUM_4;
signal  MULTS_4_6:MULT_X_SUM_4;
signal  MULTS_4_7:MULT_X_SUM_4;
signal  MULTS_4_8:MULT_X_SUM_4;
signal  MULTS_4_9:MULT_X_SUM_4;
signal  MULTS_4_10:MULT_X_SUM_4;
signal  MULTS_4_11:MULT_X_SUM_4;
signal  MULTS_4_12:MULT_X_SUM_4;
signal  MULTS_4_13:MULT_X_SUM_4;
signal  MULTS_4_14:MULT_X_SUM_4;
signal  MULTS_4_15:MULT_X_SUM_4;
signal  MULTS_4_16:MULT_X_SUM_4;
signal  MULTS_4_17:MULT_X_SUM_4;
signal  MULTS_4_18:MULT_X_SUM_4;
signal  MULTS_4_19:MULT_X_SUM_4;
signal  MULTS_4_20:MULT_X_SUM_4;
signal  MULTS_4_21:MULT_X_SUM_4;
signal  MULTS_4_22:MULT_X_SUM_4;
signal  MULTS_4_23:MULT_X_SUM_4;
signal  MULTS_4_24:MULT_X_SUM_4;
signal  MULTS_4_25:MULT_X_SUM_4;
signal  MULTS_4_26:MULT_X_SUM_4;
signal  MULTS_4_27:MULT_X_SUM_4;
signal  MULTS_4_28:MULT_X_SUM_4;
signal  MULTS_4_29:MULT_X_SUM_4;
signal  MULTS_4_30:MULT_X_SUM_4;
signal  MULTS_4_31:MULT_X_SUM_4;
signal  MULTS_4_32:MULT_X_SUM_4;
signal  MULTS_4_33:MULT_X_SUM_4;
signal  MULTS_4_34:MULT_X_SUM_4;
signal  MULTS_4_35:MULT_X_SUM_4;
signal  MULTS_4_36:MULT_X_SUM_4;
signal  MULTS_4_37:MULT_X_SUM_4;
signal  MULTS_4_38:MULT_X_SUM_4;
signal  MULTS_4_39:MULT_X_SUM_4;
signal  MULTS_4_40:MULT_X_SUM_4;
signal  MULTS_4_41:MULT_X_SUM_4;
signal  MULTS_4_42:MULT_X_SUM_4;
signal  MULTS_4_43:MULT_X_SUM_4;
signal  MULTS_4_44:MULT_X_SUM_4;
signal  MULTS_4_45:MULT_X_SUM_4;
signal  MULTS_4_46:MULT_X_SUM_4;
signal  MULTS_4_47:MULT_X_SUM_4;
signal  MULTS_4_48:MULT_X_SUM_4;
signal  MULTS_4_49:MULT_X_SUM_4;
signal  MULTS_4_50:MULT_X_SUM_4;
signal  MULTS_4_51:MULT_X_SUM_4;
signal  MULTS_4_52:MULT_X_SUM_4;
signal  MULTS_4_53:MULT_X_SUM_4;
signal  MULTS_4_54:MULT_X_SUM_4;
signal  MULTS_4_55:MULT_X_SUM_4;
signal  MULTS_4_56:MULT_X_SUM_4;
signal  MULTS_4_57:MULT_X_SUM_4;
signal  MULTS_4_58:MULT_X_SUM_4;
signal  MULTS_4_59:MULT_X_SUM_4;
signal  MULTS_4_60:MULT_X_SUM_4;
signal  MULTS_4_61:MULT_X_SUM_4;
signal  MULTS_4_62:MULT_X_SUM_4;
signal  MULTS_4_63:MULT_X_SUM_4;
signal  MULTS_4_64:MULT_X_SUM_4;
signal  MULTS_4_65:MULT_X_SUM_4;
signal  MULTS_4_66:MULT_X_SUM_4;
signal  MULTS_4_67:MULT_X_SUM_4;
signal  MULTS_4_68:MULT_X_SUM_4;
signal  MULTS_4_69:MULT_X_SUM_4;
signal  MULTS_4_70:MULT_X_SUM_4;
signal  MULTS_4_71:MULT_X_SUM_4;
signal  MULTS_4_72:MULT_X_SUM_4;
signal  MULTS_4_73:MULT_X_SUM_4;
signal  MULTS_4_74:MULT_X_SUM_4;
signal  MULTS_4_75:MULT_X_SUM_4;
signal  MULTS_4_76:MULT_X_SUM_4;
signal  MULTS_4_77:MULT_X_SUM_4;
signal  MULTS_4_78:MULT_X_SUM_4;
signal  MULTS_4_79:MULT_X_SUM_4;
signal  MULTS_4_80:MULT_X_SUM_4;
signal  MULTS_4_81:MULT_X_SUM_4;
signal  MULTS_4_82:MULT_X_SUM_4;
signal  MULTS_4_83:MULT_X_SUM_4;
signal  MULTS_4_84:MULT_X_SUM_4;
signal  MULTS_4_85:MULT_X_SUM_4;
signal  MULTS_4_86:MULT_X_SUM_4;
signal  MULTS_4_87:MULT_X_SUM_4;
signal  MULTS_4_88:MULT_X_SUM_4;
signal  MULTS_4_89:MULT_X_SUM_4;
signal  MULTS_4_90:MULT_X_SUM_4;
signal  MULTS_4_91:MULT_X_SUM_4;
signal  MULTS_4_92:MULT_X_SUM_4;
signal  MULTS_4_93:MULT_X_SUM_4;
signal  MULTS_4_94:MULT_X_SUM_4;
signal  MULTS_4_95:MULT_X_SUM_4;
signal  MULTS_4_96:MULT_X_SUM_4;
signal  MULTS_4_97:MULT_X_SUM_4;
signal  MULTS_4_98:MULT_X_SUM_4;
signal  MULTS_4_99:MULT_X_SUM_4;
signal  MULTS_4_100:MULT_X_SUM_4;
signal  MULTS_4_101:MULT_X_SUM_4;
signal  MULTS_4_102:MULT_X_SUM_4;
signal  MULTS_4_103:MULT_X_SUM_4;
signal  MULTS_4_104:MULT_X_SUM_4;
signal  MULTS_4_105:MULT_X_SUM_4;
signal  MULTS_4_106:MULT_X_SUM_4;
signal  MULTS_4_107:MULT_X_SUM_4;
signal  MULTS_4_108:MULT_X_SUM_4;
signal  MULTS_4_109:MULT_X_SUM_4;
signal  MULTS_4_110:MULT_X_SUM_4;
signal  MULTS_4_111:MULT_X_SUM_4;
signal  MULTS_4_112:MULT_X_SUM_4;
signal  MULTS_4_113:MULT_X_SUM_4;
signal  MULTS_4_114:MULT_X_SUM_4;
signal  MULTS_4_115:MULT_X_SUM_4;
signal  MULTS_4_116:MULT_X_SUM_4;
signal  MULTS_4_117:MULT_X_SUM_4;
signal  MULTS_4_118:MULT_X_SUM_4;
signal  MULTS_4_119:MULT_X_SUM_4;
signal  MULTS_4_120:MULT_X_SUM_4;
type    MULT_X_SUM_5	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_5- 1 downto 0);
signal  EN_SUM_MULT_5	: std_logic;
signal  MULTS_5_1:MULT_X_SUM_5;
signal  MULTS_5_2:MULT_X_SUM_5;
signal  MULTS_5_3:MULT_X_SUM_5;
signal  MULTS_5_4:MULT_X_SUM_5;
signal  MULTS_5_5:MULT_X_SUM_5;
signal  MULTS_5_6:MULT_X_SUM_5;
signal  MULTS_5_7:MULT_X_SUM_5;
signal  MULTS_5_8:MULT_X_SUM_5;
signal  MULTS_5_9:MULT_X_SUM_5;
signal  MULTS_5_10:MULT_X_SUM_5;
signal  MULTS_5_11:MULT_X_SUM_5;
signal  MULTS_5_12:MULT_X_SUM_5;
signal  MULTS_5_13:MULT_X_SUM_5;
signal  MULTS_5_14:MULT_X_SUM_5;
signal  MULTS_5_15:MULT_X_SUM_5;
signal  MULTS_5_16:MULT_X_SUM_5;
signal  MULTS_5_17:MULT_X_SUM_5;
signal  MULTS_5_18:MULT_X_SUM_5;
signal  MULTS_5_19:MULT_X_SUM_5;
signal  MULTS_5_20:MULT_X_SUM_5;
signal  MULTS_5_21:MULT_X_SUM_5;
signal  MULTS_5_22:MULT_X_SUM_5;
signal  MULTS_5_23:MULT_X_SUM_5;
signal  MULTS_5_24:MULT_X_SUM_5;
signal  MULTS_5_25:MULT_X_SUM_5;
signal  MULTS_5_26:MULT_X_SUM_5;
signal  MULTS_5_27:MULT_X_SUM_5;
signal  MULTS_5_28:MULT_X_SUM_5;
signal  MULTS_5_29:MULT_X_SUM_5;
signal  MULTS_5_30:MULT_X_SUM_5;
signal  MULTS_5_31:MULT_X_SUM_5;
signal  MULTS_5_32:MULT_X_SUM_5;
signal  MULTS_5_33:MULT_X_SUM_5;
signal  MULTS_5_34:MULT_X_SUM_5;
signal  MULTS_5_35:MULT_X_SUM_5;
signal  MULTS_5_36:MULT_X_SUM_5;
signal  MULTS_5_37:MULT_X_SUM_5;
signal  MULTS_5_38:MULT_X_SUM_5;
signal  MULTS_5_39:MULT_X_SUM_5;
signal  MULTS_5_40:MULT_X_SUM_5;
signal  MULTS_5_41:MULT_X_SUM_5;
signal  MULTS_5_42:MULT_X_SUM_5;
signal  MULTS_5_43:MULT_X_SUM_5;
signal  MULTS_5_44:MULT_X_SUM_5;
signal  MULTS_5_45:MULT_X_SUM_5;
signal  MULTS_5_46:MULT_X_SUM_5;
signal  MULTS_5_47:MULT_X_SUM_5;
signal  MULTS_5_48:MULT_X_SUM_5;
signal  MULTS_5_49:MULT_X_SUM_5;
signal  MULTS_5_50:MULT_X_SUM_5;
signal  MULTS_5_51:MULT_X_SUM_5;
signal  MULTS_5_52:MULT_X_SUM_5;
signal  MULTS_5_53:MULT_X_SUM_5;
signal  MULTS_5_54:MULT_X_SUM_5;
signal  MULTS_5_55:MULT_X_SUM_5;
signal  MULTS_5_56:MULT_X_SUM_5;
signal  MULTS_5_57:MULT_X_SUM_5;
signal  MULTS_5_58:MULT_X_SUM_5;
signal  MULTS_5_59:MULT_X_SUM_5;
signal  MULTS_5_60:MULT_X_SUM_5;
signal  MULTS_5_61:MULT_X_SUM_5;
signal  MULTS_5_62:MULT_X_SUM_5;
signal  MULTS_5_63:MULT_X_SUM_5;
signal  MULTS_5_64:MULT_X_SUM_5;
signal  MULTS_5_65:MULT_X_SUM_5;
signal  MULTS_5_66:MULT_X_SUM_5;
signal  MULTS_5_67:MULT_X_SUM_5;
signal  MULTS_5_68:MULT_X_SUM_5;
signal  MULTS_5_69:MULT_X_SUM_5;
signal  MULTS_5_70:MULT_X_SUM_5;
signal  MULTS_5_71:MULT_X_SUM_5;
signal  MULTS_5_72:MULT_X_SUM_5;
signal  MULTS_5_73:MULT_X_SUM_5;
signal  MULTS_5_74:MULT_X_SUM_5;
signal  MULTS_5_75:MULT_X_SUM_5;
signal  MULTS_5_76:MULT_X_SUM_5;
signal  MULTS_5_77:MULT_X_SUM_5;
signal  MULTS_5_78:MULT_X_SUM_5;
signal  MULTS_5_79:MULT_X_SUM_5;
signal  MULTS_5_80:MULT_X_SUM_5;
signal  MULTS_5_81:MULT_X_SUM_5;
signal  MULTS_5_82:MULT_X_SUM_5;
signal  MULTS_5_83:MULT_X_SUM_5;
signal  MULTS_5_84:MULT_X_SUM_5;
signal  MULTS_5_85:MULT_X_SUM_5;
signal  MULTS_5_86:MULT_X_SUM_5;
signal  MULTS_5_87:MULT_X_SUM_5;
signal  MULTS_5_88:MULT_X_SUM_5;
signal  MULTS_5_89:MULT_X_SUM_5;
signal  MULTS_5_90:MULT_X_SUM_5;
signal  MULTS_5_91:MULT_X_SUM_5;
signal  MULTS_5_92:MULT_X_SUM_5;
signal  MULTS_5_93:MULT_X_SUM_5;
signal  MULTS_5_94:MULT_X_SUM_5;
signal  MULTS_5_95:MULT_X_SUM_5;
signal  MULTS_5_96:MULT_X_SUM_5;
signal  MULTS_5_97:MULT_X_SUM_5;
signal  MULTS_5_98:MULT_X_SUM_5;
signal  MULTS_5_99:MULT_X_SUM_5;
signal  MULTS_5_100:MULT_X_SUM_5;
signal  MULTS_5_101:MULT_X_SUM_5;
signal  MULTS_5_102:MULT_X_SUM_5;
signal  MULTS_5_103:MULT_X_SUM_5;
signal  MULTS_5_104:MULT_X_SUM_5;
signal  MULTS_5_105:MULT_X_SUM_5;
signal  MULTS_5_106:MULT_X_SUM_5;
signal  MULTS_5_107:MULT_X_SUM_5;
signal  MULTS_5_108:MULT_X_SUM_5;
signal  MULTS_5_109:MULT_X_SUM_5;
signal  MULTS_5_110:MULT_X_SUM_5;
signal  MULTS_5_111:MULT_X_SUM_5;
signal  MULTS_5_112:MULT_X_SUM_5;
signal  MULTS_5_113:MULT_X_SUM_5;
signal  MULTS_5_114:MULT_X_SUM_5;
signal  MULTS_5_115:MULT_X_SUM_5;
signal  MULTS_5_116:MULT_X_SUM_5;
signal  MULTS_5_117:MULT_X_SUM_5;
signal  MULTS_5_118:MULT_X_SUM_5;
signal  MULTS_5_119:MULT_X_SUM_5;
signal  MULTS_5_120:MULT_X_SUM_5;
type    MULT_X_SUM_6	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_6- 1 downto 0);
signal  EN_SUM_MULT_6	: std_logic;
signal  MULTS_6_1:MULT_X_SUM_6;
signal  MULTS_6_2:MULT_X_SUM_6;
signal  MULTS_6_3:MULT_X_SUM_6;
signal  MULTS_6_4:MULT_X_SUM_6;
signal  MULTS_6_5:MULT_X_SUM_6;
signal  MULTS_6_6:MULT_X_SUM_6;
signal  MULTS_6_7:MULT_X_SUM_6;
signal  MULTS_6_8:MULT_X_SUM_6;
signal  MULTS_6_9:MULT_X_SUM_6;
signal  MULTS_6_10:MULT_X_SUM_6;
signal  MULTS_6_11:MULT_X_SUM_6;
signal  MULTS_6_12:MULT_X_SUM_6;
signal  MULTS_6_13:MULT_X_SUM_6;
signal  MULTS_6_14:MULT_X_SUM_6;
signal  MULTS_6_15:MULT_X_SUM_6;
signal  MULTS_6_16:MULT_X_SUM_6;
signal  MULTS_6_17:MULT_X_SUM_6;
signal  MULTS_6_18:MULT_X_SUM_6;
signal  MULTS_6_19:MULT_X_SUM_6;
signal  MULTS_6_20:MULT_X_SUM_6;
signal  MULTS_6_21:MULT_X_SUM_6;
signal  MULTS_6_22:MULT_X_SUM_6;
signal  MULTS_6_23:MULT_X_SUM_6;
signal  MULTS_6_24:MULT_X_SUM_6;
signal  MULTS_6_25:MULT_X_SUM_6;
signal  MULTS_6_26:MULT_X_SUM_6;
signal  MULTS_6_27:MULT_X_SUM_6;
signal  MULTS_6_28:MULT_X_SUM_6;
signal  MULTS_6_29:MULT_X_SUM_6;
signal  MULTS_6_30:MULT_X_SUM_6;
signal  MULTS_6_31:MULT_X_SUM_6;
signal  MULTS_6_32:MULT_X_SUM_6;
signal  MULTS_6_33:MULT_X_SUM_6;
signal  MULTS_6_34:MULT_X_SUM_6;
signal  MULTS_6_35:MULT_X_SUM_6;
signal  MULTS_6_36:MULT_X_SUM_6;
signal  MULTS_6_37:MULT_X_SUM_6;
signal  MULTS_6_38:MULT_X_SUM_6;
signal  MULTS_6_39:MULT_X_SUM_6;
signal  MULTS_6_40:MULT_X_SUM_6;
signal  MULTS_6_41:MULT_X_SUM_6;
signal  MULTS_6_42:MULT_X_SUM_6;
signal  MULTS_6_43:MULT_X_SUM_6;
signal  MULTS_6_44:MULT_X_SUM_6;
signal  MULTS_6_45:MULT_X_SUM_6;
signal  MULTS_6_46:MULT_X_SUM_6;
signal  MULTS_6_47:MULT_X_SUM_6;
signal  MULTS_6_48:MULT_X_SUM_6;
signal  MULTS_6_49:MULT_X_SUM_6;
signal  MULTS_6_50:MULT_X_SUM_6;
signal  MULTS_6_51:MULT_X_SUM_6;
signal  MULTS_6_52:MULT_X_SUM_6;
signal  MULTS_6_53:MULT_X_SUM_6;
signal  MULTS_6_54:MULT_X_SUM_6;
signal  MULTS_6_55:MULT_X_SUM_6;
signal  MULTS_6_56:MULT_X_SUM_6;
signal  MULTS_6_57:MULT_X_SUM_6;
signal  MULTS_6_58:MULT_X_SUM_6;
signal  MULTS_6_59:MULT_X_SUM_6;
signal  MULTS_6_60:MULT_X_SUM_6;
signal  MULTS_6_61:MULT_X_SUM_6;
signal  MULTS_6_62:MULT_X_SUM_6;
signal  MULTS_6_63:MULT_X_SUM_6;
signal  MULTS_6_64:MULT_X_SUM_6;
signal  MULTS_6_65:MULT_X_SUM_6;
signal  MULTS_6_66:MULT_X_SUM_6;
signal  MULTS_6_67:MULT_X_SUM_6;
signal  MULTS_6_68:MULT_X_SUM_6;
signal  MULTS_6_69:MULT_X_SUM_6;
signal  MULTS_6_70:MULT_X_SUM_6;
signal  MULTS_6_71:MULT_X_SUM_6;
signal  MULTS_6_72:MULT_X_SUM_6;
signal  MULTS_6_73:MULT_X_SUM_6;
signal  MULTS_6_74:MULT_X_SUM_6;
signal  MULTS_6_75:MULT_X_SUM_6;
signal  MULTS_6_76:MULT_X_SUM_6;
signal  MULTS_6_77:MULT_X_SUM_6;
signal  MULTS_6_78:MULT_X_SUM_6;
signal  MULTS_6_79:MULT_X_SUM_6;
signal  MULTS_6_80:MULT_X_SUM_6;
signal  MULTS_6_81:MULT_X_SUM_6;
signal  MULTS_6_82:MULT_X_SUM_6;
signal  MULTS_6_83:MULT_X_SUM_6;
signal  MULTS_6_84:MULT_X_SUM_6;
signal  MULTS_6_85:MULT_X_SUM_6;
signal  MULTS_6_86:MULT_X_SUM_6;
signal  MULTS_6_87:MULT_X_SUM_6;
signal  MULTS_6_88:MULT_X_SUM_6;
signal  MULTS_6_89:MULT_X_SUM_6;
signal  MULTS_6_90:MULT_X_SUM_6;
signal  MULTS_6_91:MULT_X_SUM_6;
signal  MULTS_6_92:MULT_X_SUM_6;
signal  MULTS_6_93:MULT_X_SUM_6;
signal  MULTS_6_94:MULT_X_SUM_6;
signal  MULTS_6_95:MULT_X_SUM_6;
signal  MULTS_6_96:MULT_X_SUM_6;
signal  MULTS_6_97:MULT_X_SUM_6;
signal  MULTS_6_98:MULT_X_SUM_6;
signal  MULTS_6_99:MULT_X_SUM_6;
signal  MULTS_6_100:MULT_X_SUM_6;
signal  MULTS_6_101:MULT_X_SUM_6;
signal  MULTS_6_102:MULT_X_SUM_6;
signal  MULTS_6_103:MULT_X_SUM_6;
signal  MULTS_6_104:MULT_X_SUM_6;
signal  MULTS_6_105:MULT_X_SUM_6;
signal  MULTS_6_106:MULT_X_SUM_6;
signal  MULTS_6_107:MULT_X_SUM_6;
signal  MULTS_6_108:MULT_X_SUM_6;
signal  MULTS_6_109:MULT_X_SUM_6;
signal  MULTS_6_110:MULT_X_SUM_6;
signal  MULTS_6_111:MULT_X_SUM_6;
signal  MULTS_6_112:MULT_X_SUM_6;
signal  MULTS_6_113:MULT_X_SUM_6;
signal  MULTS_6_114:MULT_X_SUM_6;
signal  MULTS_6_115:MULT_X_SUM_6;
signal  MULTS_6_116:MULT_X_SUM_6;
signal  MULTS_6_117:MULT_X_SUM_6;
signal  MULTS_6_118:MULT_X_SUM_6;
signal  MULTS_6_119:MULT_X_SUM_6;
signal  MULTS_6_120:MULT_X_SUM_6;
type    MULT_X_SUM_7	is array (0 to FEATURE_MAPS-1 ) of signed(MULT_SUM_SIZE_7- 1 downto 0);
signal  EN_SUM_MULT_7	: std_logic;
signal  MULTS_7_1:MULT_X_SUM_7;
signal  MULTS_7_2:MULT_X_SUM_7;
signal  MULTS_7_3:MULT_X_SUM_7;
signal  MULTS_7_4:MULT_X_SUM_7;
signal  MULTS_7_5:MULT_X_SUM_7;
signal  MULTS_7_6:MULT_X_SUM_7;
signal  MULTS_7_7:MULT_X_SUM_7;
signal  MULTS_7_8:MULT_X_SUM_7;
signal  MULTS_7_9:MULT_X_SUM_7;
signal  MULTS_7_10:MULT_X_SUM_7;
signal  MULTS_7_11:MULT_X_SUM_7;
signal  MULTS_7_12:MULT_X_SUM_7;
signal  MULTS_7_13:MULT_X_SUM_7;
signal  MULTS_7_14:MULT_X_SUM_7;
signal  MULTS_7_15:MULT_X_SUM_7;
signal  MULTS_7_16:MULT_X_SUM_7;
signal  MULTS_7_17:MULT_X_SUM_7;
signal  MULTS_7_18:MULT_X_SUM_7;
signal  MULTS_7_19:MULT_X_SUM_7;
signal  MULTS_7_20:MULT_X_SUM_7;
signal  MULTS_7_21:MULT_X_SUM_7;
signal  MULTS_7_22:MULT_X_SUM_7;
signal  MULTS_7_23:MULT_X_SUM_7;
signal  MULTS_7_24:MULT_X_SUM_7;
signal  MULTS_7_25:MULT_X_SUM_7;
signal  MULTS_7_26:MULT_X_SUM_7;
signal  MULTS_7_27:MULT_X_SUM_7;
signal  MULTS_7_28:MULT_X_SUM_7;
signal  MULTS_7_29:MULT_X_SUM_7;
signal  MULTS_7_30:MULT_X_SUM_7;
signal  MULTS_7_31:MULT_X_SUM_7;
signal  MULTS_7_32:MULT_X_SUM_7;
signal  MULTS_7_33:MULT_X_SUM_7;
signal  MULTS_7_34:MULT_X_SUM_7;
signal  MULTS_7_35:MULT_X_SUM_7;
signal  MULTS_7_36:MULT_X_SUM_7;
signal  MULTS_7_37:MULT_X_SUM_7;
signal  MULTS_7_38:MULT_X_SUM_7;
signal  MULTS_7_39:MULT_X_SUM_7;
signal  MULTS_7_40:MULT_X_SUM_7;
signal  MULTS_7_41:MULT_X_SUM_7;
signal  MULTS_7_42:MULT_X_SUM_7;
signal  MULTS_7_43:MULT_X_SUM_7;
signal  MULTS_7_44:MULT_X_SUM_7;
signal  MULTS_7_45:MULT_X_SUM_7;
signal  MULTS_7_46:MULT_X_SUM_7;
signal  MULTS_7_47:MULT_X_SUM_7;
signal  MULTS_7_48:MULT_X_SUM_7;
signal  MULTS_7_49:MULT_X_SUM_7;
signal  MULTS_7_50:MULT_X_SUM_7;
signal  MULTS_7_51:MULT_X_SUM_7;
signal  MULTS_7_52:MULT_X_SUM_7;
signal  MULTS_7_53:MULT_X_SUM_7;
signal  MULTS_7_54:MULT_X_SUM_7;
signal  MULTS_7_55:MULT_X_SUM_7;
signal  MULTS_7_56:MULT_X_SUM_7;
signal  MULTS_7_57:MULT_X_SUM_7;
signal  MULTS_7_58:MULT_X_SUM_7;
signal  MULTS_7_59:MULT_X_SUM_7;
signal  MULTS_7_60:MULT_X_SUM_7;
signal  MULTS_7_61:MULT_X_SUM_7;
signal  MULTS_7_62:MULT_X_SUM_7;
signal  MULTS_7_63:MULT_X_SUM_7;
signal  MULTS_7_64:MULT_X_SUM_7;
signal  MULTS_7_65:MULT_X_SUM_7;
signal  MULTS_7_66:MULT_X_SUM_7;
signal  MULTS_7_67:MULT_X_SUM_7;
signal  MULTS_7_68:MULT_X_SUM_7;
signal  MULTS_7_69:MULT_X_SUM_7;
signal  MULTS_7_70:MULT_X_SUM_7;
signal  MULTS_7_71:MULT_X_SUM_7;
signal  MULTS_7_72:MULT_X_SUM_7;
signal  MULTS_7_73:MULT_X_SUM_7;
signal  MULTS_7_74:MULT_X_SUM_7;
signal  MULTS_7_75:MULT_X_SUM_7;
signal  MULTS_7_76:MULT_X_SUM_7;
signal  MULTS_7_77:MULT_X_SUM_7;
signal  MULTS_7_78:MULT_X_SUM_7;
signal  MULTS_7_79:MULT_X_SUM_7;
signal  MULTS_7_80:MULT_X_SUM_7;
signal  MULTS_7_81:MULT_X_SUM_7;
signal  MULTS_7_82:MULT_X_SUM_7;
signal  MULTS_7_83:MULT_X_SUM_7;
signal  MULTS_7_84:MULT_X_SUM_7;
signal  MULTS_7_85:MULT_X_SUM_7;
signal  MULTS_7_86:MULT_X_SUM_7;
signal  MULTS_7_87:MULT_X_SUM_7;
signal  MULTS_7_88:MULT_X_SUM_7;
signal  MULTS_7_89:MULT_X_SUM_7;
signal  MULTS_7_90:MULT_X_SUM_7;
signal  MULTS_7_91:MULT_X_SUM_7;
signal  MULTS_7_92:MULT_X_SUM_7;
signal  MULTS_7_93:MULT_X_SUM_7;
signal  MULTS_7_94:MULT_X_SUM_7;
signal  MULTS_7_95:MULT_X_SUM_7;
signal  MULTS_7_96:MULT_X_SUM_7;
signal  MULTS_7_97:MULT_X_SUM_7;
signal  MULTS_7_98:MULT_X_SUM_7;
signal  MULTS_7_99:MULT_X_SUM_7;
signal  MULTS_7_100:MULT_X_SUM_7;
signal  MULTS_7_101:MULT_X_SUM_7;
signal  MULTS_7_102:MULT_X_SUM_7;
signal  MULTS_7_103:MULT_X_SUM_7;
signal  MULTS_7_104:MULT_X_SUM_7;
signal  MULTS_7_105:MULT_X_SUM_7;
signal  MULTS_7_106:MULT_X_SUM_7;
signal  MULTS_7_107:MULT_X_SUM_7;
signal  MULTS_7_108:MULT_X_SUM_7;
signal  MULTS_7_109:MULT_X_SUM_7;
signal  MULTS_7_110:MULT_X_SUM_7;
signal  MULTS_7_111:MULT_X_SUM_7;
signal  MULTS_7_112:MULT_X_SUM_7;
signal  MULTS_7_113:MULT_X_SUM_7;
signal  MULTS_7_114:MULT_X_SUM_7;
signal  MULTS_7_115:MULT_X_SUM_7;
signal  MULTS_7_116:MULT_X_SUM_7;
signal  MULTS_7_117:MULT_X_SUM_7;
signal  MULTS_7_118:MULT_X_SUM_7;
signal  MULTS_7_119:MULT_X_SUM_7;
signal  MULTS_7_120:MULT_X_SUM_7;


-------------------------------------- OUTPUT FROM LOWER COMPONENT SIGNALS--------------------------------------------------
signal DOUT_1_8          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_2_8          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_3_8          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_4_8          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_5_8          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_6_8          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_7_8          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_8_8          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_9_8          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_10_8          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal EN_STREAM_OUT_8	 : std_logic;
signal VALID_OUT_8       : std_logic;

--------------------------------------------- FILTER HARDCODED CONSTANTS -WEIGHTS START--------------------------------

constant FMAP_1_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_11_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_12_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_13_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_14_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_15_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_16_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_17_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_18_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_19_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_20_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_21_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_22_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_23_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_24_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_25_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_26_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_27_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_28_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_29_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_30_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_31_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_32_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_33_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_34_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_35_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_36_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_37_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_38_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_39_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_40_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_41_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_42_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_43_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_44_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_45_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_46_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_47_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_48_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_49_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_50_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_51_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_52_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_53_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_54_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_55_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_56_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_57_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_58_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_59_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_60_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_61_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_62_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_63_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_64_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_65_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_66_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_67_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_68_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_69_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_70_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_71_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_72_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_73_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_74_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_75_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_76_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_77_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_78_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_79_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_80_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_81_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_82_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_83_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_84_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";

constant BIAS_VAL_1: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_2: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_3: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_4: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_5: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_6: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_7: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_8: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_9: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_10: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_11: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_12: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_13: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_14: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_15: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_16: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_17: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_18: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_19: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_20: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_21: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_22: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_23: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_24: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_25: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_26: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_27: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_28: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_29: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_30: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_31: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_32: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_33: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_34: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_35: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_36: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_37: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_38: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_39: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_40: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_41: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_42: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_43: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_44: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_45: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_46: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_47: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_48: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_49: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_50: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_51: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_52: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_53: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_54: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_55: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_56: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_57: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_58: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_59: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_60: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_61: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_62: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_63: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_64: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_65: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_66: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_67: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_68: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_69: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_70: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_71: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_72: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_73: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_74: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_75: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_76: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_77: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_78: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_79: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_80: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_81: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_82: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_83: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_84: signed (BIASES_SIZE-1 downto 0):="01";


---------------------------------- MAP NEXT LAYER - COMPONENTS START----------------------------------
COMPONENT FC_LAYER_8
    port(	CLK,RST			:IN std_logic;
		DIN_1_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_2_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_3_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_4_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_5_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_6_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_7_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_8_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_9_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_10_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_11_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_12_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_13_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_14_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_15_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_16_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_17_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_18_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_19_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_20_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_21_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_22_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_23_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_24_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_25_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_26_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_27_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_28_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_29_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_30_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_31_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_32_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_33_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_34_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_35_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_36_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_37_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_38_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_39_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_40_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_41_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_42_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_43_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_44_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_45_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_46_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_47_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_48_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_49_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_50_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_51_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_52_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_53_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_54_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_55_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_56_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_57_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_58_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_59_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_60_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_61_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_62_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_63_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_64_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_65_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_66_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_67_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_68_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_69_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_70_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_71_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_72_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_73_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_74_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_75_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_76_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_77_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_78_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_79_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_80_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_81_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_82_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_83_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_84_8		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		EN_STREAM_OUT_8	:OUT std_logic;
		VALID_OUT_8		:OUT std_logic;
		DOUT_1_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_2_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_3_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_4_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_5_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_6_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_7_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_8_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_9_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_10_8        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		EN_STREAM		:IN std_logic;
		EN_LOC_STREAM_8	:IN std_logic
      			);
END COMPONENT FC_LAYER_8;

begin

FC_LYR_8 : FC_LAYER_8 
          port map(
          CLK                 => CLK,
          RST                 => RST,
          DIN_1_8             => DOUT_BUF_1_7,
          DIN_2_8             => DOUT_BUF_2_7,
          DIN_3_8             => DOUT_BUF_3_7,
          DIN_4_8             => DOUT_BUF_4_7,
          DIN_5_8             => DOUT_BUF_5_7,
          DIN_6_8             => DOUT_BUF_6_7,
          DIN_7_8             => DOUT_BUF_7_7,
          DIN_8_8             => DOUT_BUF_8_7,
          DIN_9_8             => DOUT_BUF_9_7,
          DIN_10_8             => DOUT_BUF_10_7,
          DIN_11_8             => DOUT_BUF_11_7,
          DIN_12_8             => DOUT_BUF_12_7,
          DIN_13_8             => DOUT_BUF_13_7,
          DIN_14_8             => DOUT_BUF_14_7,
          DIN_15_8             => DOUT_BUF_15_7,
          DIN_16_8             => DOUT_BUF_16_7,
          DIN_17_8             => DOUT_BUF_17_7,
          DIN_18_8             => DOUT_BUF_18_7,
          DIN_19_8             => DOUT_BUF_19_7,
          DIN_20_8             => DOUT_BUF_20_7,
          DIN_21_8             => DOUT_BUF_21_7,
          DIN_22_8             => DOUT_BUF_22_7,
          DIN_23_8             => DOUT_BUF_23_7,
          DIN_24_8             => DOUT_BUF_24_7,
          DIN_25_8             => DOUT_BUF_25_7,
          DIN_26_8             => DOUT_BUF_26_7,
          DIN_27_8             => DOUT_BUF_27_7,
          DIN_28_8             => DOUT_BUF_28_7,
          DIN_29_8             => DOUT_BUF_29_7,
          DIN_30_8             => DOUT_BUF_30_7,
          DIN_31_8             => DOUT_BUF_31_7,
          DIN_32_8             => DOUT_BUF_32_7,
          DIN_33_8             => DOUT_BUF_33_7,
          DIN_34_8             => DOUT_BUF_34_7,
          DIN_35_8             => DOUT_BUF_35_7,
          DIN_36_8             => DOUT_BUF_36_7,
          DIN_37_8             => DOUT_BUF_37_7,
          DIN_38_8             => DOUT_BUF_38_7,
          DIN_39_8             => DOUT_BUF_39_7,
          DIN_40_8             => DOUT_BUF_40_7,
          DIN_41_8             => DOUT_BUF_41_7,
          DIN_42_8             => DOUT_BUF_42_7,
          DIN_43_8             => DOUT_BUF_43_7,
          DIN_44_8             => DOUT_BUF_44_7,
          DIN_45_8             => DOUT_BUF_45_7,
          DIN_46_8             => DOUT_BUF_46_7,
          DIN_47_8             => DOUT_BUF_47_7,
          DIN_48_8             => DOUT_BUF_48_7,
          DIN_49_8             => DOUT_BUF_49_7,
          DIN_50_8             => DOUT_BUF_50_7,
          DIN_51_8             => DOUT_BUF_51_7,
          DIN_52_8             => DOUT_BUF_52_7,
          DIN_53_8             => DOUT_BUF_53_7,
          DIN_54_8             => DOUT_BUF_54_7,
          DIN_55_8             => DOUT_BUF_55_7,
          DIN_56_8             => DOUT_BUF_56_7,
          DIN_57_8             => DOUT_BUF_57_7,
          DIN_58_8             => DOUT_BUF_58_7,
          DIN_59_8             => DOUT_BUF_59_7,
          DIN_60_8             => DOUT_BUF_60_7,
          DIN_61_8             => DOUT_BUF_61_7,
          DIN_62_8             => DOUT_BUF_62_7,
          DIN_63_8             => DOUT_BUF_63_7,
          DIN_64_8             => DOUT_BUF_64_7,
          DIN_65_8             => DOUT_BUF_65_7,
          DIN_66_8             => DOUT_BUF_66_7,
          DIN_67_8             => DOUT_BUF_67_7,
          DIN_68_8             => DOUT_BUF_68_7,
          DIN_69_8             => DOUT_BUF_69_7,
          DIN_70_8             => DOUT_BUF_70_7,
          DIN_71_8             => DOUT_BUF_71_7,
          DIN_72_8             => DOUT_BUF_72_7,
          DIN_73_8             => DOUT_BUF_73_7,
          DIN_74_8             => DOUT_BUF_74_7,
          DIN_75_8             => DOUT_BUF_75_7,
          DIN_76_8             => DOUT_BUF_76_7,
          DIN_77_8             => DOUT_BUF_77_7,
          DIN_78_8             => DOUT_BUF_78_7,
          DIN_79_8             => DOUT_BUF_79_7,
          DIN_80_8             => DOUT_BUF_80_7,
          DIN_81_8             => DOUT_BUF_81_7,
          DIN_82_8             => DOUT_BUF_82_7,
          DIN_83_8             => DOUT_BUF_83_7,
          DIN_84_8             => DOUT_BUF_84_7,
          DOUT_1_8            => DOUT_1_8,
          DOUT_2_8            => DOUT_2_8,
          DOUT_3_8            => DOUT_3_8,
          DOUT_4_8            => DOUT_4_8,
          DOUT_5_8            => DOUT_5_8,
          DOUT_6_8            => DOUT_6_8,
          DOUT_7_8            => DOUT_7_8,
          DOUT_8_8            => DOUT_8_8,
          DOUT_9_8            => DOUT_9_8,
          DOUT_10_8            => DOUT_10_8,
          VALID_OUT_8         => VALID_OUT_8,
          EN_STREAM_OUT_8     => EN_STREAM_OUT_8,
          EN_LOC_STREAM_8     => EN_NXT_LYR_7,
          EN_STREAM           => EN_STREAM
                );

----------------------------------------------- MAP NEXT LAYER - COMPONENTS END----------------------------------------------------



-------------------------------------------------------- ARCHITECTURE BEGIN--------------------------------------------------------

LAYER_7: process(CLK)


begin
------------------------------------------------ RESET AND PROCESS TOP START ------------------------------------------------------
if rising_edge(CLK) then
  if RST = '1' then
	-------------------FIXED SIGNALS RESET------------------------
    PIXEL_COUNT<=0;VALID_NXTLYR_PIX<=0;OUT_PIXEL_COUNT<=0;
    EN_NXT_LYR_7<='0';FRST_TIM_EN_7<='0';INTERNAL_RST<='0';
    Enable_MULT<='0';Enable_ADDER<='0';Enable_ReLU<='0';Enable_BIAS<='0';
    PADDING_count<=0;ROW_COUNT<=0;SIG_STRIDE<=STRIDE;COUNT_PIX<=0;

-------------------DYNAMIC SIGNALS RESET------------------------
    DOUT_BUF_1_7<=(others => '0');BIAS_1<=(others => '0');ReLU_1<=(others => '0');
    DOUT_BUF_2_7<=(others => '0');BIAS_2<=(others => '0');ReLU_2<=(others => '0');
    DOUT_BUF_3_7<=(others => '0');BIAS_3<=(others => '0');ReLU_3<=(others => '0');
    DOUT_BUF_4_7<=(others => '0');BIAS_4<=(others => '0');ReLU_4<=(others => '0');
    DOUT_BUF_5_7<=(others => '0');BIAS_5<=(others => '0');ReLU_5<=(others => '0');
    DOUT_BUF_6_7<=(others => '0');BIAS_6<=(others => '0');ReLU_6<=(others => '0');
    DOUT_BUF_7_7<=(others => '0');BIAS_7<=(others => '0');ReLU_7<=(others => '0');
    DOUT_BUF_8_7<=(others => '0');BIAS_8<=(others => '0');ReLU_8<=(others => '0');
    DOUT_BUF_9_7<=(others => '0');BIAS_9<=(others => '0');ReLU_9<=(others => '0');
    DOUT_BUF_10_7<=(others => '0');BIAS_10<=(others => '0');ReLU_10<=(others => '0');
    DOUT_BUF_11_7<=(others => '0');BIAS_11<=(others => '0');ReLU_11<=(others => '0');
    DOUT_BUF_12_7<=(others => '0');BIAS_12<=(others => '0');ReLU_12<=(others => '0');
    DOUT_BUF_13_7<=(others => '0');BIAS_13<=(others => '0');ReLU_13<=(others => '0');
    DOUT_BUF_14_7<=(others => '0');BIAS_14<=(others => '0');ReLU_14<=(others => '0');
    DOUT_BUF_15_7<=(others => '0');BIAS_15<=(others => '0');ReLU_15<=(others => '0');
    DOUT_BUF_16_7<=(others => '0');BIAS_16<=(others => '0');ReLU_16<=(others => '0');
    DOUT_BUF_17_7<=(others => '0');BIAS_17<=(others => '0');ReLU_17<=(others => '0');
    DOUT_BUF_18_7<=(others => '0');BIAS_18<=(others => '0');ReLU_18<=(others => '0');
    DOUT_BUF_19_7<=(others => '0');BIAS_19<=(others => '0');ReLU_19<=(others => '0');
    DOUT_BUF_20_7<=(others => '0');BIAS_20<=(others => '0');ReLU_20<=(others => '0');
    DOUT_BUF_21_7<=(others => '0');BIAS_21<=(others => '0');ReLU_21<=(others => '0');
    DOUT_BUF_22_7<=(others => '0');BIAS_22<=(others => '0');ReLU_22<=(others => '0');
    DOUT_BUF_23_7<=(others => '0');BIAS_23<=(others => '0');ReLU_23<=(others => '0');
    DOUT_BUF_24_7<=(others => '0');BIAS_24<=(others => '0');ReLU_24<=(others => '0');
    DOUT_BUF_25_7<=(others => '0');BIAS_25<=(others => '0');ReLU_25<=(others => '0');
    DOUT_BUF_26_7<=(others => '0');BIAS_26<=(others => '0');ReLU_26<=(others => '0');
    DOUT_BUF_27_7<=(others => '0');BIAS_27<=(others => '0');ReLU_27<=(others => '0');
    DOUT_BUF_28_7<=(others => '0');BIAS_28<=(others => '0');ReLU_28<=(others => '0');
    DOUT_BUF_29_7<=(others => '0');BIAS_29<=(others => '0');ReLU_29<=(others => '0');
    DOUT_BUF_30_7<=(others => '0');BIAS_30<=(others => '0');ReLU_30<=(others => '0');
    DOUT_BUF_31_7<=(others => '0');BIAS_31<=(others => '0');ReLU_31<=(others => '0');
    DOUT_BUF_32_7<=(others => '0');BIAS_32<=(others => '0');ReLU_32<=(others => '0');
    DOUT_BUF_33_7<=(others => '0');BIAS_33<=(others => '0');ReLU_33<=(others => '0');
    DOUT_BUF_34_7<=(others => '0');BIAS_34<=(others => '0');ReLU_34<=(others => '0');
    DOUT_BUF_35_7<=(others => '0');BIAS_35<=(others => '0');ReLU_35<=(others => '0');
    DOUT_BUF_36_7<=(others => '0');BIAS_36<=(others => '0');ReLU_36<=(others => '0');
    DOUT_BUF_37_7<=(others => '0');BIAS_37<=(others => '0');ReLU_37<=(others => '0');
    DOUT_BUF_38_7<=(others => '0');BIAS_38<=(others => '0');ReLU_38<=(others => '0');
    DOUT_BUF_39_7<=(others => '0');BIAS_39<=(others => '0');ReLU_39<=(others => '0');
    DOUT_BUF_40_7<=(others => '0');BIAS_40<=(others => '0');ReLU_40<=(others => '0');
    DOUT_BUF_41_7<=(others => '0');BIAS_41<=(others => '0');ReLU_41<=(others => '0');
    DOUT_BUF_42_7<=(others => '0');BIAS_42<=(others => '0');ReLU_42<=(others => '0');
    DOUT_BUF_43_7<=(others => '0');BIAS_43<=(others => '0');ReLU_43<=(others => '0');
    DOUT_BUF_44_7<=(others => '0');BIAS_44<=(others => '0');ReLU_44<=(others => '0');
    DOUT_BUF_45_7<=(others => '0');BIAS_45<=(others => '0');ReLU_45<=(others => '0');
    DOUT_BUF_46_7<=(others => '0');BIAS_46<=(others => '0');ReLU_46<=(others => '0');
    DOUT_BUF_47_7<=(others => '0');BIAS_47<=(others => '0');ReLU_47<=(others => '0');
    DOUT_BUF_48_7<=(others => '0');BIAS_48<=(others => '0');ReLU_48<=(others => '0');
    DOUT_BUF_49_7<=(others => '0');BIAS_49<=(others => '0');ReLU_49<=(others => '0');
    DOUT_BUF_50_7<=(others => '0');BIAS_50<=(others => '0');ReLU_50<=(others => '0');
    DOUT_BUF_51_7<=(others => '0');BIAS_51<=(others => '0');ReLU_51<=(others => '0');
    DOUT_BUF_52_7<=(others => '0');BIAS_52<=(others => '0');ReLU_52<=(others => '0');
    DOUT_BUF_53_7<=(others => '0');BIAS_53<=(others => '0');ReLU_53<=(others => '0');
    DOUT_BUF_54_7<=(others => '0');BIAS_54<=(others => '0');ReLU_54<=(others => '0');
    DOUT_BUF_55_7<=(others => '0');BIAS_55<=(others => '0');ReLU_55<=(others => '0');
    DOUT_BUF_56_7<=(others => '0');BIAS_56<=(others => '0');ReLU_56<=(others => '0');
    DOUT_BUF_57_7<=(others => '0');BIAS_57<=(others => '0');ReLU_57<=(others => '0');
    DOUT_BUF_58_7<=(others => '0');BIAS_58<=(others => '0');ReLU_58<=(others => '0');
    DOUT_BUF_59_7<=(others => '0');BIAS_59<=(others => '0');ReLU_59<=(others => '0');
    DOUT_BUF_60_7<=(others => '0');BIAS_60<=(others => '0');ReLU_60<=(others => '0');
    DOUT_BUF_61_7<=(others => '0');BIAS_61<=(others => '0');ReLU_61<=(others => '0');
    DOUT_BUF_62_7<=(others => '0');BIAS_62<=(others => '0');ReLU_62<=(others => '0');
    DOUT_BUF_63_7<=(others => '0');BIAS_63<=(others => '0');ReLU_63<=(others => '0');
    DOUT_BUF_64_7<=(others => '0');BIAS_64<=(others => '0');ReLU_64<=(others => '0');
    DOUT_BUF_65_7<=(others => '0');BIAS_65<=(others => '0');ReLU_65<=(others => '0');
    DOUT_BUF_66_7<=(others => '0');BIAS_66<=(others => '0');ReLU_66<=(others => '0');
    DOUT_BUF_67_7<=(others => '0');BIAS_67<=(others => '0');ReLU_67<=(others => '0');
    DOUT_BUF_68_7<=(others => '0');BIAS_68<=(others => '0');ReLU_68<=(others => '0');
    DOUT_BUF_69_7<=(others => '0');BIAS_69<=(others => '0');ReLU_69<=(others => '0');
    DOUT_BUF_70_7<=(others => '0');BIAS_70<=(others => '0');ReLU_70<=(others => '0');
    DOUT_BUF_71_7<=(others => '0');BIAS_71<=(others => '0');ReLU_71<=(others => '0');
    DOUT_BUF_72_7<=(others => '0');BIAS_72<=(others => '0');ReLU_72<=(others => '0');
    DOUT_BUF_73_7<=(others => '0');BIAS_73<=(others => '0');ReLU_73<=(others => '0');
    DOUT_BUF_74_7<=(others => '0');BIAS_74<=(others => '0');ReLU_74<=(others => '0');
    DOUT_BUF_75_7<=(others => '0');BIAS_75<=(others => '0');ReLU_75<=(others => '0');
    DOUT_BUF_76_7<=(others => '0');BIAS_76<=(others => '0');ReLU_76<=(others => '0');
    DOUT_BUF_77_7<=(others => '0');BIAS_77<=(others => '0');ReLU_77<=(others => '0');
    DOUT_BUF_78_7<=(others => '0');BIAS_78<=(others => '0');ReLU_78<=(others => '0');
    DOUT_BUF_79_7<=(others => '0');BIAS_79<=(others => '0');ReLU_79<=(others => '0');
    DOUT_BUF_80_7<=(others => '0');BIAS_80<=(others => '0');ReLU_80<=(others => '0');
    DOUT_BUF_81_7<=(others => '0');BIAS_81<=(others => '0');ReLU_81<=(others => '0');
    DOUT_BUF_82_7<=(others => '0');BIAS_82<=(others => '0');ReLU_82<=(others => '0');
    DOUT_BUF_83_7<=(others => '0');BIAS_83<=(others => '0');ReLU_83<=(others => '0');
    DOUT_BUF_84_7<=(others => '0');BIAS_84<=(others => '0');ReLU_84<=(others => '0');

    SUM_PIXELS_1<=(others=>'0');MULT_1<=((others=> (others=>'0')));
    SUM_PIXELS_2<=(others=>'0');MULT_2<=((others=> (others=>'0')));
    SUM_PIXELS_3<=(others=>'0');MULT_3<=((others=> (others=>'0')));
    SUM_PIXELS_4<=(others=>'0');MULT_4<=((others=> (others=>'0')));
    SUM_PIXELS_5<=(others=>'0');MULT_5<=((others=> (others=>'0')));
    SUM_PIXELS_6<=(others=>'0');MULT_6<=((others=> (others=>'0')));
    SUM_PIXELS_7<=(others=>'0');MULT_7<=((others=> (others=>'0')));
    SUM_PIXELS_8<=(others=>'0');MULT_8<=((others=> (others=>'0')));
    SUM_PIXELS_9<=(others=>'0');MULT_9<=((others=> (others=>'0')));
    SUM_PIXELS_10<=(others=>'0');MULT_10<=((others=> (others=>'0')));
    SUM_PIXELS_11<=(others=>'0');MULT_11<=((others=> (others=>'0')));
    SUM_PIXELS_12<=(others=>'0');MULT_12<=((others=> (others=>'0')));
    SUM_PIXELS_13<=(others=>'0');MULT_13<=((others=> (others=>'0')));
    SUM_PIXELS_14<=(others=>'0');MULT_14<=((others=> (others=>'0')));
    SUM_PIXELS_15<=(others=>'0');MULT_15<=((others=> (others=>'0')));
    SUM_PIXELS_16<=(others=>'0');MULT_16<=((others=> (others=>'0')));
    SUM_PIXELS_17<=(others=>'0');MULT_17<=((others=> (others=>'0')));
    SUM_PIXELS_18<=(others=>'0');MULT_18<=((others=> (others=>'0')));
    SUM_PIXELS_19<=(others=>'0');MULT_19<=((others=> (others=>'0')));
    SUM_PIXELS_20<=(others=>'0');MULT_20<=((others=> (others=>'0')));
    SUM_PIXELS_21<=(others=>'0');MULT_21<=((others=> (others=>'0')));
    SUM_PIXELS_22<=(others=>'0');MULT_22<=((others=> (others=>'0')));
    SUM_PIXELS_23<=(others=>'0');MULT_23<=((others=> (others=>'0')));
    SUM_PIXELS_24<=(others=>'0');MULT_24<=((others=> (others=>'0')));
    SUM_PIXELS_25<=(others=>'0');MULT_25<=((others=> (others=>'0')));
    SUM_PIXELS_26<=(others=>'0');MULT_26<=((others=> (others=>'0')));
    SUM_PIXELS_27<=(others=>'0');MULT_27<=((others=> (others=>'0')));
    SUM_PIXELS_28<=(others=>'0');MULT_28<=((others=> (others=>'0')));
    SUM_PIXELS_29<=(others=>'0');MULT_29<=((others=> (others=>'0')));
    SUM_PIXELS_30<=(others=>'0');MULT_30<=((others=> (others=>'0')));
    SUM_PIXELS_31<=(others=>'0');MULT_31<=((others=> (others=>'0')));
    SUM_PIXELS_32<=(others=>'0');MULT_32<=((others=> (others=>'0')));
    SUM_PIXELS_33<=(others=>'0');MULT_33<=((others=> (others=>'0')));
    SUM_PIXELS_34<=(others=>'0');MULT_34<=((others=> (others=>'0')));
    SUM_PIXELS_35<=(others=>'0');MULT_35<=((others=> (others=>'0')));
    SUM_PIXELS_36<=(others=>'0');MULT_36<=((others=> (others=>'0')));
    SUM_PIXELS_37<=(others=>'0');MULT_37<=((others=> (others=>'0')));
    SUM_PIXELS_38<=(others=>'0');MULT_38<=((others=> (others=>'0')));
    SUM_PIXELS_39<=(others=>'0');MULT_39<=((others=> (others=>'0')));
    SUM_PIXELS_40<=(others=>'0');MULT_40<=((others=> (others=>'0')));
    SUM_PIXELS_41<=(others=>'0');MULT_41<=((others=> (others=>'0')));
    SUM_PIXELS_42<=(others=>'0');MULT_42<=((others=> (others=>'0')));
    SUM_PIXELS_43<=(others=>'0');MULT_43<=((others=> (others=>'0')));
    SUM_PIXELS_44<=(others=>'0');MULT_44<=((others=> (others=>'0')));
    SUM_PIXELS_45<=(others=>'0');MULT_45<=((others=> (others=>'0')));
    SUM_PIXELS_46<=(others=>'0');MULT_46<=((others=> (others=>'0')));
    SUM_PIXELS_47<=(others=>'0');MULT_47<=((others=> (others=>'0')));
    SUM_PIXELS_48<=(others=>'0');MULT_48<=((others=> (others=>'0')));
    SUM_PIXELS_49<=(others=>'0');MULT_49<=((others=> (others=>'0')));
    SUM_PIXELS_50<=(others=>'0');MULT_50<=((others=> (others=>'0')));
    SUM_PIXELS_51<=(others=>'0');MULT_51<=((others=> (others=>'0')));
    SUM_PIXELS_52<=(others=>'0');MULT_52<=((others=> (others=>'0')));
    SUM_PIXELS_53<=(others=>'0');MULT_53<=((others=> (others=>'0')));
    SUM_PIXELS_54<=(others=>'0');MULT_54<=((others=> (others=>'0')));
    SUM_PIXELS_55<=(others=>'0');MULT_55<=((others=> (others=>'0')));
    SUM_PIXELS_56<=(others=>'0');MULT_56<=((others=> (others=>'0')));
    SUM_PIXELS_57<=(others=>'0');MULT_57<=((others=> (others=>'0')));
    SUM_PIXELS_58<=(others=>'0');MULT_58<=((others=> (others=>'0')));
    SUM_PIXELS_59<=(others=>'0');MULT_59<=((others=> (others=>'0')));
    SUM_PIXELS_60<=(others=>'0');MULT_60<=((others=> (others=>'0')));
    SUM_PIXELS_61<=(others=>'0');MULT_61<=((others=> (others=>'0')));
    SUM_PIXELS_62<=(others=>'0');MULT_62<=((others=> (others=>'0')));
    SUM_PIXELS_63<=(others=>'0');MULT_63<=((others=> (others=>'0')));
    SUM_PIXELS_64<=(others=>'0');MULT_64<=((others=> (others=>'0')));
    SUM_PIXELS_65<=(others=>'0');MULT_65<=((others=> (others=>'0')));
    SUM_PIXELS_66<=(others=>'0');MULT_66<=((others=> (others=>'0')));
    SUM_PIXELS_67<=(others=>'0');MULT_67<=((others=> (others=>'0')));
    SUM_PIXELS_68<=(others=>'0');MULT_68<=((others=> (others=>'0')));
    SUM_PIXELS_69<=(others=>'0');MULT_69<=((others=> (others=>'0')));
    SUM_PIXELS_70<=(others=>'0');MULT_70<=((others=> (others=>'0')));
    SUM_PIXELS_71<=(others=>'0');MULT_71<=((others=> (others=>'0')));
    SUM_PIXELS_72<=(others=>'0');MULT_72<=((others=> (others=>'0')));
    SUM_PIXELS_73<=(others=>'0');MULT_73<=((others=> (others=>'0')));
    SUM_PIXELS_74<=(others=>'0');MULT_74<=((others=> (others=>'0')));
    SUM_PIXELS_75<=(others=>'0');MULT_75<=((others=> (others=>'0')));
    SUM_PIXELS_76<=(others=>'0');MULT_76<=((others=> (others=>'0')));
    SUM_PIXELS_77<=(others=>'0');MULT_77<=((others=> (others=>'0')));
    SUM_PIXELS_78<=(others=>'0');MULT_78<=((others=> (others=>'0')));
    SUM_PIXELS_79<=(others=>'0');MULT_79<=((others=> (others=>'0')));
    SUM_PIXELS_80<=(others=>'0');MULT_80<=((others=> (others=>'0')));
    SUM_PIXELS_81<=(others=>'0');MULT_81<=((others=> (others=>'0')));
    SUM_PIXELS_82<=(others=>'0');MULT_82<=((others=> (others=>'0')));
    SUM_PIXELS_83<=(others=>'0');MULT_83<=((others=> (others=>'0')));
    SUM_PIXELS_84<=(others=>'0');MULT_84<=((others=> (others=>'0')));
    SUM_PIXELS_85<=(others=>'0');MULT_85<=((others=> (others=>'0')));
    SUM_PIXELS_86<=(others=>'0');MULT_86<=((others=> (others=>'0')));
    SUM_PIXELS_87<=(others=>'0');MULT_87<=((others=> (others=>'0')));
    SUM_PIXELS_88<=(others=>'0');MULT_88<=((others=> (others=>'0')));
    SUM_PIXELS_89<=(others=>'0');MULT_89<=((others=> (others=>'0')));
    SUM_PIXELS_90<=(others=>'0');MULT_90<=((others=> (others=>'0')));
    SUM_PIXELS_91<=(others=>'0');MULT_91<=((others=> (others=>'0')));
    SUM_PIXELS_92<=(others=>'0');MULT_92<=((others=> (others=>'0')));
    SUM_PIXELS_93<=(others=>'0');MULT_93<=((others=> (others=>'0')));
    SUM_PIXELS_94<=(others=>'0');MULT_94<=((others=> (others=>'0')));
    SUM_PIXELS_95<=(others=>'0');MULT_95<=((others=> (others=>'0')));
    SUM_PIXELS_96<=(others=>'0');MULT_96<=((others=> (others=>'0')));
    SUM_PIXELS_97<=(others=>'0');MULT_97<=((others=> (others=>'0')));
    SUM_PIXELS_98<=(others=>'0');MULT_98<=((others=> (others=>'0')));
    SUM_PIXELS_99<=(others=>'0');MULT_99<=((others=> (others=>'0')));
    SUM_PIXELS_100<=(others=>'0');MULT_100<=((others=> (others=>'0')));
    SUM_PIXELS_101<=(others=>'0');MULT_101<=((others=> (others=>'0')));
    SUM_PIXELS_102<=(others=>'0');MULT_102<=((others=> (others=>'0')));
    SUM_PIXELS_103<=(others=>'0');MULT_103<=((others=> (others=>'0')));
    SUM_PIXELS_104<=(others=>'0');MULT_104<=((others=> (others=>'0')));
    SUM_PIXELS_105<=(others=>'0');MULT_105<=((others=> (others=>'0')));
    SUM_PIXELS_106<=(others=>'0');MULT_106<=((others=> (others=>'0')));
    SUM_PIXELS_107<=(others=>'0');MULT_107<=((others=> (others=>'0')));
    SUM_PIXELS_108<=(others=>'0');MULT_108<=((others=> (others=>'0')));
    SUM_PIXELS_109<=(others=>'0');MULT_109<=((others=> (others=>'0')));
    SUM_PIXELS_110<=(others=>'0');MULT_110<=((others=> (others=>'0')));
    SUM_PIXELS_111<=(others=>'0');MULT_111<=((others=> (others=>'0')));
    SUM_PIXELS_112<=(others=>'0');MULT_112<=((others=> (others=>'0')));
    SUM_PIXELS_113<=(others=>'0');MULT_113<=((others=> (others=>'0')));
    SUM_PIXELS_114<=(others=>'0');MULT_114<=((others=> (others=>'0')));
    SUM_PIXELS_115<=(others=>'0');MULT_115<=((others=> (others=>'0')));
    SUM_PIXELS_116<=(others=>'0');MULT_116<=((others=> (others=>'0')));
    SUM_PIXELS_117<=(others=>'0');MULT_117<=((others=> (others=>'0')));
    SUM_PIXELS_118<=(others=>'0');MULT_118<=((others=> (others=>'0')));
    SUM_PIXELS_119<=(others=>'0');MULT_119<=((others=> (others=>'0')));
    SUM_PIXELS_120<=(others=>'0');MULT_120<=((others=> (others=>'0')));

    EN_SUM_MULT_1<='0';
    MULTS_1_1<=((others=> (others=>'0')));
    MULTS_1_2<=((others=> (others=>'0')));
    MULTS_1_3<=((others=> (others=>'0')));
    MULTS_1_4<=((others=> (others=>'0')));
    MULTS_1_5<=((others=> (others=>'0')));
    MULTS_1_6<=((others=> (others=>'0')));
    MULTS_1_7<=((others=> (others=>'0')));
    MULTS_1_8<=((others=> (others=>'0')));
    MULTS_1_9<=((others=> (others=>'0')));
    MULTS_1_10<=((others=> (others=>'0')));
    MULTS_1_11<=((others=> (others=>'0')));
    MULTS_1_12<=((others=> (others=>'0')));
    MULTS_1_13<=((others=> (others=>'0')));
    MULTS_1_14<=((others=> (others=>'0')));
    MULTS_1_15<=((others=> (others=>'0')));
    MULTS_1_16<=((others=> (others=>'0')));
    MULTS_1_17<=((others=> (others=>'0')));
    MULTS_1_18<=((others=> (others=>'0')));
    MULTS_1_19<=((others=> (others=>'0')));
    MULTS_1_20<=((others=> (others=>'0')));
    MULTS_1_21<=((others=> (others=>'0')));
    MULTS_1_22<=((others=> (others=>'0')));
    MULTS_1_23<=((others=> (others=>'0')));
    MULTS_1_24<=((others=> (others=>'0')));
    MULTS_1_25<=((others=> (others=>'0')));
    MULTS_1_26<=((others=> (others=>'0')));
    MULTS_1_27<=((others=> (others=>'0')));
    MULTS_1_28<=((others=> (others=>'0')));
    MULTS_1_29<=((others=> (others=>'0')));
    MULTS_1_30<=((others=> (others=>'0')));
    MULTS_1_31<=((others=> (others=>'0')));
    MULTS_1_32<=((others=> (others=>'0')));
    MULTS_1_33<=((others=> (others=>'0')));
    MULTS_1_34<=((others=> (others=>'0')));
    MULTS_1_35<=((others=> (others=>'0')));
    MULTS_1_36<=((others=> (others=>'0')));
    MULTS_1_37<=((others=> (others=>'0')));
    MULTS_1_38<=((others=> (others=>'0')));
    MULTS_1_39<=((others=> (others=>'0')));
    MULTS_1_40<=((others=> (others=>'0')));
    MULTS_1_41<=((others=> (others=>'0')));
    MULTS_1_42<=((others=> (others=>'0')));
    MULTS_1_43<=((others=> (others=>'0')));
    MULTS_1_44<=((others=> (others=>'0')));
    MULTS_1_45<=((others=> (others=>'0')));
    MULTS_1_46<=((others=> (others=>'0')));
    MULTS_1_47<=((others=> (others=>'0')));
    MULTS_1_48<=((others=> (others=>'0')));
    MULTS_1_49<=((others=> (others=>'0')));
    MULTS_1_50<=((others=> (others=>'0')));
    MULTS_1_51<=((others=> (others=>'0')));
    MULTS_1_52<=((others=> (others=>'0')));
    MULTS_1_53<=((others=> (others=>'0')));
    MULTS_1_54<=((others=> (others=>'0')));
    MULTS_1_55<=((others=> (others=>'0')));
    MULTS_1_56<=((others=> (others=>'0')));
    MULTS_1_57<=((others=> (others=>'0')));
    MULTS_1_58<=((others=> (others=>'0')));
    MULTS_1_59<=((others=> (others=>'0')));
    MULTS_1_60<=((others=> (others=>'0')));
    MULTS_1_61<=((others=> (others=>'0')));
    MULTS_1_62<=((others=> (others=>'0')));
    MULTS_1_63<=((others=> (others=>'0')));
    MULTS_1_64<=((others=> (others=>'0')));
    MULTS_1_65<=((others=> (others=>'0')));
    MULTS_1_66<=((others=> (others=>'0')));
    MULTS_1_67<=((others=> (others=>'0')));
    MULTS_1_68<=((others=> (others=>'0')));
    MULTS_1_69<=((others=> (others=>'0')));
    MULTS_1_70<=((others=> (others=>'0')));
    MULTS_1_71<=((others=> (others=>'0')));
    MULTS_1_72<=((others=> (others=>'0')));
    MULTS_1_73<=((others=> (others=>'0')));
    MULTS_1_74<=((others=> (others=>'0')));
    MULTS_1_75<=((others=> (others=>'0')));
    MULTS_1_76<=((others=> (others=>'0')));
    MULTS_1_77<=((others=> (others=>'0')));
    MULTS_1_78<=((others=> (others=>'0')));
    MULTS_1_79<=((others=> (others=>'0')));
    MULTS_1_80<=((others=> (others=>'0')));
    MULTS_1_81<=((others=> (others=>'0')));
    MULTS_1_82<=((others=> (others=>'0')));
    MULTS_1_83<=((others=> (others=>'0')));
    MULTS_1_84<=((others=> (others=>'0')));
    MULTS_1_85<=((others=> (others=>'0')));
    MULTS_1_86<=((others=> (others=>'0')));
    MULTS_1_87<=((others=> (others=>'0')));
    MULTS_1_88<=((others=> (others=>'0')));
    MULTS_1_89<=((others=> (others=>'0')));
    MULTS_1_90<=((others=> (others=>'0')));
    MULTS_1_91<=((others=> (others=>'0')));
    MULTS_1_92<=((others=> (others=>'0')));
    MULTS_1_93<=((others=> (others=>'0')));
    MULTS_1_94<=((others=> (others=>'0')));
    MULTS_1_95<=((others=> (others=>'0')));
    MULTS_1_96<=((others=> (others=>'0')));
    MULTS_1_97<=((others=> (others=>'0')));
    MULTS_1_98<=((others=> (others=>'0')));
    MULTS_1_99<=((others=> (others=>'0')));
    MULTS_1_100<=((others=> (others=>'0')));
    MULTS_1_101<=((others=> (others=>'0')));
    MULTS_1_102<=((others=> (others=>'0')));
    MULTS_1_103<=((others=> (others=>'0')));
    MULTS_1_104<=((others=> (others=>'0')));
    MULTS_1_105<=((others=> (others=>'0')));
    MULTS_1_106<=((others=> (others=>'0')));
    MULTS_1_107<=((others=> (others=>'0')));
    MULTS_1_108<=((others=> (others=>'0')));
    MULTS_1_109<=((others=> (others=>'0')));
    MULTS_1_110<=((others=> (others=>'0')));
    MULTS_1_111<=((others=> (others=>'0')));
    MULTS_1_112<=((others=> (others=>'0')));
    MULTS_1_113<=((others=> (others=>'0')));
    MULTS_1_114<=((others=> (others=>'0')));
    MULTS_1_115<=((others=> (others=>'0')));
    MULTS_1_116<=((others=> (others=>'0')));
    MULTS_1_117<=((others=> (others=>'0')));
    MULTS_1_118<=((others=> (others=>'0')));
    MULTS_1_119<=((others=> (others=>'0')));
    MULTS_1_120<=((others=> (others=>'0')));
    EN_SUM_MULT_2<='0';
    MULTS_2_1<=((others=> (others=>'0')));
    MULTS_2_2<=((others=> (others=>'0')));
    MULTS_2_3<=((others=> (others=>'0')));
    MULTS_2_4<=((others=> (others=>'0')));
    MULTS_2_5<=((others=> (others=>'0')));
    MULTS_2_6<=((others=> (others=>'0')));
    MULTS_2_7<=((others=> (others=>'0')));
    MULTS_2_8<=((others=> (others=>'0')));
    MULTS_2_9<=((others=> (others=>'0')));
    MULTS_2_10<=((others=> (others=>'0')));
    MULTS_2_11<=((others=> (others=>'0')));
    MULTS_2_12<=((others=> (others=>'0')));
    MULTS_2_13<=((others=> (others=>'0')));
    MULTS_2_14<=((others=> (others=>'0')));
    MULTS_2_15<=((others=> (others=>'0')));
    MULTS_2_16<=((others=> (others=>'0')));
    MULTS_2_17<=((others=> (others=>'0')));
    MULTS_2_18<=((others=> (others=>'0')));
    MULTS_2_19<=((others=> (others=>'0')));
    MULTS_2_20<=((others=> (others=>'0')));
    MULTS_2_21<=((others=> (others=>'0')));
    MULTS_2_22<=((others=> (others=>'0')));
    MULTS_2_23<=((others=> (others=>'0')));
    MULTS_2_24<=((others=> (others=>'0')));
    MULTS_2_25<=((others=> (others=>'0')));
    MULTS_2_26<=((others=> (others=>'0')));
    MULTS_2_27<=((others=> (others=>'0')));
    MULTS_2_28<=((others=> (others=>'0')));
    MULTS_2_29<=((others=> (others=>'0')));
    MULTS_2_30<=((others=> (others=>'0')));
    MULTS_2_31<=((others=> (others=>'0')));
    MULTS_2_32<=((others=> (others=>'0')));
    MULTS_2_33<=((others=> (others=>'0')));
    MULTS_2_34<=((others=> (others=>'0')));
    MULTS_2_35<=((others=> (others=>'0')));
    MULTS_2_36<=((others=> (others=>'0')));
    MULTS_2_37<=((others=> (others=>'0')));
    MULTS_2_38<=((others=> (others=>'0')));
    MULTS_2_39<=((others=> (others=>'0')));
    MULTS_2_40<=((others=> (others=>'0')));
    MULTS_2_41<=((others=> (others=>'0')));
    MULTS_2_42<=((others=> (others=>'0')));
    MULTS_2_43<=((others=> (others=>'0')));
    MULTS_2_44<=((others=> (others=>'0')));
    MULTS_2_45<=((others=> (others=>'0')));
    MULTS_2_46<=((others=> (others=>'0')));
    MULTS_2_47<=((others=> (others=>'0')));
    MULTS_2_48<=((others=> (others=>'0')));
    MULTS_2_49<=((others=> (others=>'0')));
    MULTS_2_50<=((others=> (others=>'0')));
    MULTS_2_51<=((others=> (others=>'0')));
    MULTS_2_52<=((others=> (others=>'0')));
    MULTS_2_53<=((others=> (others=>'0')));
    MULTS_2_54<=((others=> (others=>'0')));
    MULTS_2_55<=((others=> (others=>'0')));
    MULTS_2_56<=((others=> (others=>'0')));
    MULTS_2_57<=((others=> (others=>'0')));
    MULTS_2_58<=((others=> (others=>'0')));
    MULTS_2_59<=((others=> (others=>'0')));
    MULTS_2_60<=((others=> (others=>'0')));
    MULTS_2_61<=((others=> (others=>'0')));
    MULTS_2_62<=((others=> (others=>'0')));
    MULTS_2_63<=((others=> (others=>'0')));
    MULTS_2_64<=((others=> (others=>'0')));
    MULTS_2_65<=((others=> (others=>'0')));
    MULTS_2_66<=((others=> (others=>'0')));
    MULTS_2_67<=((others=> (others=>'0')));
    MULTS_2_68<=((others=> (others=>'0')));
    MULTS_2_69<=((others=> (others=>'0')));
    MULTS_2_70<=((others=> (others=>'0')));
    MULTS_2_71<=((others=> (others=>'0')));
    MULTS_2_72<=((others=> (others=>'0')));
    MULTS_2_73<=((others=> (others=>'0')));
    MULTS_2_74<=((others=> (others=>'0')));
    MULTS_2_75<=((others=> (others=>'0')));
    MULTS_2_76<=((others=> (others=>'0')));
    MULTS_2_77<=((others=> (others=>'0')));
    MULTS_2_78<=((others=> (others=>'0')));
    MULTS_2_79<=((others=> (others=>'0')));
    MULTS_2_80<=((others=> (others=>'0')));
    MULTS_2_81<=((others=> (others=>'0')));
    MULTS_2_82<=((others=> (others=>'0')));
    MULTS_2_83<=((others=> (others=>'0')));
    MULTS_2_84<=((others=> (others=>'0')));
    MULTS_2_85<=((others=> (others=>'0')));
    MULTS_2_86<=((others=> (others=>'0')));
    MULTS_2_87<=((others=> (others=>'0')));
    MULTS_2_88<=((others=> (others=>'0')));
    MULTS_2_89<=((others=> (others=>'0')));
    MULTS_2_90<=((others=> (others=>'0')));
    MULTS_2_91<=((others=> (others=>'0')));
    MULTS_2_92<=((others=> (others=>'0')));
    MULTS_2_93<=((others=> (others=>'0')));
    MULTS_2_94<=((others=> (others=>'0')));
    MULTS_2_95<=((others=> (others=>'0')));
    MULTS_2_96<=((others=> (others=>'0')));
    MULTS_2_97<=((others=> (others=>'0')));
    MULTS_2_98<=((others=> (others=>'0')));
    MULTS_2_99<=((others=> (others=>'0')));
    MULTS_2_100<=((others=> (others=>'0')));
    MULTS_2_101<=((others=> (others=>'0')));
    MULTS_2_102<=((others=> (others=>'0')));
    MULTS_2_103<=((others=> (others=>'0')));
    MULTS_2_104<=((others=> (others=>'0')));
    MULTS_2_105<=((others=> (others=>'0')));
    MULTS_2_106<=((others=> (others=>'0')));
    MULTS_2_107<=((others=> (others=>'0')));
    MULTS_2_108<=((others=> (others=>'0')));
    MULTS_2_109<=((others=> (others=>'0')));
    MULTS_2_110<=((others=> (others=>'0')));
    MULTS_2_111<=((others=> (others=>'0')));
    MULTS_2_112<=((others=> (others=>'0')));
    MULTS_2_113<=((others=> (others=>'0')));
    MULTS_2_114<=((others=> (others=>'0')));
    MULTS_2_115<=((others=> (others=>'0')));
    MULTS_2_116<=((others=> (others=>'0')));
    MULTS_2_117<=((others=> (others=>'0')));
    MULTS_2_118<=((others=> (others=>'0')));
    MULTS_2_119<=((others=> (others=>'0')));
    MULTS_2_120<=((others=> (others=>'0')));
    EN_SUM_MULT_3<='0';
    MULTS_3_1<=((others=> (others=>'0')));
    MULTS_3_2<=((others=> (others=>'0')));
    MULTS_3_3<=((others=> (others=>'0')));
    MULTS_3_4<=((others=> (others=>'0')));
    MULTS_3_5<=((others=> (others=>'0')));
    MULTS_3_6<=((others=> (others=>'0')));
    MULTS_3_7<=((others=> (others=>'0')));
    MULTS_3_8<=((others=> (others=>'0')));
    MULTS_3_9<=((others=> (others=>'0')));
    MULTS_3_10<=((others=> (others=>'0')));
    MULTS_3_11<=((others=> (others=>'0')));
    MULTS_3_12<=((others=> (others=>'0')));
    MULTS_3_13<=((others=> (others=>'0')));
    MULTS_3_14<=((others=> (others=>'0')));
    MULTS_3_15<=((others=> (others=>'0')));
    MULTS_3_16<=((others=> (others=>'0')));
    MULTS_3_17<=((others=> (others=>'0')));
    MULTS_3_18<=((others=> (others=>'0')));
    MULTS_3_19<=((others=> (others=>'0')));
    MULTS_3_20<=((others=> (others=>'0')));
    MULTS_3_21<=((others=> (others=>'0')));
    MULTS_3_22<=((others=> (others=>'0')));
    MULTS_3_23<=((others=> (others=>'0')));
    MULTS_3_24<=((others=> (others=>'0')));
    MULTS_3_25<=((others=> (others=>'0')));
    MULTS_3_26<=((others=> (others=>'0')));
    MULTS_3_27<=((others=> (others=>'0')));
    MULTS_3_28<=((others=> (others=>'0')));
    MULTS_3_29<=((others=> (others=>'0')));
    MULTS_3_30<=((others=> (others=>'0')));
    MULTS_3_31<=((others=> (others=>'0')));
    MULTS_3_32<=((others=> (others=>'0')));
    MULTS_3_33<=((others=> (others=>'0')));
    MULTS_3_34<=((others=> (others=>'0')));
    MULTS_3_35<=((others=> (others=>'0')));
    MULTS_3_36<=((others=> (others=>'0')));
    MULTS_3_37<=((others=> (others=>'0')));
    MULTS_3_38<=((others=> (others=>'0')));
    MULTS_3_39<=((others=> (others=>'0')));
    MULTS_3_40<=((others=> (others=>'0')));
    MULTS_3_41<=((others=> (others=>'0')));
    MULTS_3_42<=((others=> (others=>'0')));
    MULTS_3_43<=((others=> (others=>'0')));
    MULTS_3_44<=((others=> (others=>'0')));
    MULTS_3_45<=((others=> (others=>'0')));
    MULTS_3_46<=((others=> (others=>'0')));
    MULTS_3_47<=((others=> (others=>'0')));
    MULTS_3_48<=((others=> (others=>'0')));
    MULTS_3_49<=((others=> (others=>'0')));
    MULTS_3_50<=((others=> (others=>'0')));
    MULTS_3_51<=((others=> (others=>'0')));
    MULTS_3_52<=((others=> (others=>'0')));
    MULTS_3_53<=((others=> (others=>'0')));
    MULTS_3_54<=((others=> (others=>'0')));
    MULTS_3_55<=((others=> (others=>'0')));
    MULTS_3_56<=((others=> (others=>'0')));
    MULTS_3_57<=((others=> (others=>'0')));
    MULTS_3_58<=((others=> (others=>'0')));
    MULTS_3_59<=((others=> (others=>'0')));
    MULTS_3_60<=((others=> (others=>'0')));
    MULTS_3_61<=((others=> (others=>'0')));
    MULTS_3_62<=((others=> (others=>'0')));
    MULTS_3_63<=((others=> (others=>'0')));
    MULTS_3_64<=((others=> (others=>'0')));
    MULTS_3_65<=((others=> (others=>'0')));
    MULTS_3_66<=((others=> (others=>'0')));
    MULTS_3_67<=((others=> (others=>'0')));
    MULTS_3_68<=((others=> (others=>'0')));
    MULTS_3_69<=((others=> (others=>'0')));
    MULTS_3_70<=((others=> (others=>'0')));
    MULTS_3_71<=((others=> (others=>'0')));
    MULTS_3_72<=((others=> (others=>'0')));
    MULTS_3_73<=((others=> (others=>'0')));
    MULTS_3_74<=((others=> (others=>'0')));
    MULTS_3_75<=((others=> (others=>'0')));
    MULTS_3_76<=((others=> (others=>'0')));
    MULTS_3_77<=((others=> (others=>'0')));
    MULTS_3_78<=((others=> (others=>'0')));
    MULTS_3_79<=((others=> (others=>'0')));
    MULTS_3_80<=((others=> (others=>'0')));
    MULTS_3_81<=((others=> (others=>'0')));
    MULTS_3_82<=((others=> (others=>'0')));
    MULTS_3_83<=((others=> (others=>'0')));
    MULTS_3_84<=((others=> (others=>'0')));
    MULTS_3_85<=((others=> (others=>'0')));
    MULTS_3_86<=((others=> (others=>'0')));
    MULTS_3_87<=((others=> (others=>'0')));
    MULTS_3_88<=((others=> (others=>'0')));
    MULTS_3_89<=((others=> (others=>'0')));
    MULTS_3_90<=((others=> (others=>'0')));
    MULTS_3_91<=((others=> (others=>'0')));
    MULTS_3_92<=((others=> (others=>'0')));
    MULTS_3_93<=((others=> (others=>'0')));
    MULTS_3_94<=((others=> (others=>'0')));
    MULTS_3_95<=((others=> (others=>'0')));
    MULTS_3_96<=((others=> (others=>'0')));
    MULTS_3_97<=((others=> (others=>'0')));
    MULTS_3_98<=((others=> (others=>'0')));
    MULTS_3_99<=((others=> (others=>'0')));
    MULTS_3_100<=((others=> (others=>'0')));
    MULTS_3_101<=((others=> (others=>'0')));
    MULTS_3_102<=((others=> (others=>'0')));
    MULTS_3_103<=((others=> (others=>'0')));
    MULTS_3_104<=((others=> (others=>'0')));
    MULTS_3_105<=((others=> (others=>'0')));
    MULTS_3_106<=((others=> (others=>'0')));
    MULTS_3_107<=((others=> (others=>'0')));
    MULTS_3_108<=((others=> (others=>'0')));
    MULTS_3_109<=((others=> (others=>'0')));
    MULTS_3_110<=((others=> (others=>'0')));
    MULTS_3_111<=((others=> (others=>'0')));
    MULTS_3_112<=((others=> (others=>'0')));
    MULTS_3_113<=((others=> (others=>'0')));
    MULTS_3_114<=((others=> (others=>'0')));
    MULTS_3_115<=((others=> (others=>'0')));
    MULTS_3_116<=((others=> (others=>'0')));
    MULTS_3_117<=((others=> (others=>'0')));
    MULTS_3_118<=((others=> (others=>'0')));
    MULTS_3_119<=((others=> (others=>'0')));
    MULTS_3_120<=((others=> (others=>'0')));
    EN_SUM_MULT_4<='0';
    MULTS_4_1<=((others=> (others=>'0')));
    MULTS_4_2<=((others=> (others=>'0')));
    MULTS_4_3<=((others=> (others=>'0')));
    MULTS_4_4<=((others=> (others=>'0')));
    MULTS_4_5<=((others=> (others=>'0')));
    MULTS_4_6<=((others=> (others=>'0')));
    MULTS_4_7<=((others=> (others=>'0')));
    MULTS_4_8<=((others=> (others=>'0')));
    MULTS_4_9<=((others=> (others=>'0')));
    MULTS_4_10<=((others=> (others=>'0')));
    MULTS_4_11<=((others=> (others=>'0')));
    MULTS_4_12<=((others=> (others=>'0')));
    MULTS_4_13<=((others=> (others=>'0')));
    MULTS_4_14<=((others=> (others=>'0')));
    MULTS_4_15<=((others=> (others=>'0')));
    MULTS_4_16<=((others=> (others=>'0')));
    MULTS_4_17<=((others=> (others=>'0')));
    MULTS_4_18<=((others=> (others=>'0')));
    MULTS_4_19<=((others=> (others=>'0')));
    MULTS_4_20<=((others=> (others=>'0')));
    MULTS_4_21<=((others=> (others=>'0')));
    MULTS_4_22<=((others=> (others=>'0')));
    MULTS_4_23<=((others=> (others=>'0')));
    MULTS_4_24<=((others=> (others=>'0')));
    MULTS_4_25<=((others=> (others=>'0')));
    MULTS_4_26<=((others=> (others=>'0')));
    MULTS_4_27<=((others=> (others=>'0')));
    MULTS_4_28<=((others=> (others=>'0')));
    MULTS_4_29<=((others=> (others=>'0')));
    MULTS_4_30<=((others=> (others=>'0')));
    MULTS_4_31<=((others=> (others=>'0')));
    MULTS_4_32<=((others=> (others=>'0')));
    MULTS_4_33<=((others=> (others=>'0')));
    MULTS_4_34<=((others=> (others=>'0')));
    MULTS_4_35<=((others=> (others=>'0')));
    MULTS_4_36<=((others=> (others=>'0')));
    MULTS_4_37<=((others=> (others=>'0')));
    MULTS_4_38<=((others=> (others=>'0')));
    MULTS_4_39<=((others=> (others=>'0')));
    MULTS_4_40<=((others=> (others=>'0')));
    MULTS_4_41<=((others=> (others=>'0')));
    MULTS_4_42<=((others=> (others=>'0')));
    MULTS_4_43<=((others=> (others=>'0')));
    MULTS_4_44<=((others=> (others=>'0')));
    MULTS_4_45<=((others=> (others=>'0')));
    MULTS_4_46<=((others=> (others=>'0')));
    MULTS_4_47<=((others=> (others=>'0')));
    MULTS_4_48<=((others=> (others=>'0')));
    MULTS_4_49<=((others=> (others=>'0')));
    MULTS_4_50<=((others=> (others=>'0')));
    MULTS_4_51<=((others=> (others=>'0')));
    MULTS_4_52<=((others=> (others=>'0')));
    MULTS_4_53<=((others=> (others=>'0')));
    MULTS_4_54<=((others=> (others=>'0')));
    MULTS_4_55<=((others=> (others=>'0')));
    MULTS_4_56<=((others=> (others=>'0')));
    MULTS_4_57<=((others=> (others=>'0')));
    MULTS_4_58<=((others=> (others=>'0')));
    MULTS_4_59<=((others=> (others=>'0')));
    MULTS_4_60<=((others=> (others=>'0')));
    MULTS_4_61<=((others=> (others=>'0')));
    MULTS_4_62<=((others=> (others=>'0')));
    MULTS_4_63<=((others=> (others=>'0')));
    MULTS_4_64<=((others=> (others=>'0')));
    MULTS_4_65<=((others=> (others=>'0')));
    MULTS_4_66<=((others=> (others=>'0')));
    MULTS_4_67<=((others=> (others=>'0')));
    MULTS_4_68<=((others=> (others=>'0')));
    MULTS_4_69<=((others=> (others=>'0')));
    MULTS_4_70<=((others=> (others=>'0')));
    MULTS_4_71<=((others=> (others=>'0')));
    MULTS_4_72<=((others=> (others=>'0')));
    MULTS_4_73<=((others=> (others=>'0')));
    MULTS_4_74<=((others=> (others=>'0')));
    MULTS_4_75<=((others=> (others=>'0')));
    MULTS_4_76<=((others=> (others=>'0')));
    MULTS_4_77<=((others=> (others=>'0')));
    MULTS_4_78<=((others=> (others=>'0')));
    MULTS_4_79<=((others=> (others=>'0')));
    MULTS_4_80<=((others=> (others=>'0')));
    MULTS_4_81<=((others=> (others=>'0')));
    MULTS_4_82<=((others=> (others=>'0')));
    MULTS_4_83<=((others=> (others=>'0')));
    MULTS_4_84<=((others=> (others=>'0')));
    MULTS_4_85<=((others=> (others=>'0')));
    MULTS_4_86<=((others=> (others=>'0')));
    MULTS_4_87<=((others=> (others=>'0')));
    MULTS_4_88<=((others=> (others=>'0')));
    MULTS_4_89<=((others=> (others=>'0')));
    MULTS_4_90<=((others=> (others=>'0')));
    MULTS_4_91<=((others=> (others=>'0')));
    MULTS_4_92<=((others=> (others=>'0')));
    MULTS_4_93<=((others=> (others=>'0')));
    MULTS_4_94<=((others=> (others=>'0')));
    MULTS_4_95<=((others=> (others=>'0')));
    MULTS_4_96<=((others=> (others=>'0')));
    MULTS_4_97<=((others=> (others=>'0')));
    MULTS_4_98<=((others=> (others=>'0')));
    MULTS_4_99<=((others=> (others=>'0')));
    MULTS_4_100<=((others=> (others=>'0')));
    MULTS_4_101<=((others=> (others=>'0')));
    MULTS_4_102<=((others=> (others=>'0')));
    MULTS_4_103<=((others=> (others=>'0')));
    MULTS_4_104<=((others=> (others=>'0')));
    MULTS_4_105<=((others=> (others=>'0')));
    MULTS_4_106<=((others=> (others=>'0')));
    MULTS_4_107<=((others=> (others=>'0')));
    MULTS_4_108<=((others=> (others=>'0')));
    MULTS_4_109<=((others=> (others=>'0')));
    MULTS_4_110<=((others=> (others=>'0')));
    MULTS_4_111<=((others=> (others=>'0')));
    MULTS_4_112<=((others=> (others=>'0')));
    MULTS_4_113<=((others=> (others=>'0')));
    MULTS_4_114<=((others=> (others=>'0')));
    MULTS_4_115<=((others=> (others=>'0')));
    MULTS_4_116<=((others=> (others=>'0')));
    MULTS_4_117<=((others=> (others=>'0')));
    MULTS_4_118<=((others=> (others=>'0')));
    MULTS_4_119<=((others=> (others=>'0')));
    MULTS_4_120<=((others=> (others=>'0')));
    EN_SUM_MULT_5<='0';
    MULTS_5_1<=((others=> (others=>'0')));
    MULTS_5_2<=((others=> (others=>'0')));
    MULTS_5_3<=((others=> (others=>'0')));
    MULTS_5_4<=((others=> (others=>'0')));
    MULTS_5_5<=((others=> (others=>'0')));
    MULTS_5_6<=((others=> (others=>'0')));
    MULTS_5_7<=((others=> (others=>'0')));
    MULTS_5_8<=((others=> (others=>'0')));
    MULTS_5_9<=((others=> (others=>'0')));
    MULTS_5_10<=((others=> (others=>'0')));
    MULTS_5_11<=((others=> (others=>'0')));
    MULTS_5_12<=((others=> (others=>'0')));
    MULTS_5_13<=((others=> (others=>'0')));
    MULTS_5_14<=((others=> (others=>'0')));
    MULTS_5_15<=((others=> (others=>'0')));
    MULTS_5_16<=((others=> (others=>'0')));
    MULTS_5_17<=((others=> (others=>'0')));
    MULTS_5_18<=((others=> (others=>'0')));
    MULTS_5_19<=((others=> (others=>'0')));
    MULTS_5_20<=((others=> (others=>'0')));
    MULTS_5_21<=((others=> (others=>'0')));
    MULTS_5_22<=((others=> (others=>'0')));
    MULTS_5_23<=((others=> (others=>'0')));
    MULTS_5_24<=((others=> (others=>'0')));
    MULTS_5_25<=((others=> (others=>'0')));
    MULTS_5_26<=((others=> (others=>'0')));
    MULTS_5_27<=((others=> (others=>'0')));
    MULTS_5_28<=((others=> (others=>'0')));
    MULTS_5_29<=((others=> (others=>'0')));
    MULTS_5_30<=((others=> (others=>'0')));
    MULTS_5_31<=((others=> (others=>'0')));
    MULTS_5_32<=((others=> (others=>'0')));
    MULTS_5_33<=((others=> (others=>'0')));
    MULTS_5_34<=((others=> (others=>'0')));
    MULTS_5_35<=((others=> (others=>'0')));
    MULTS_5_36<=((others=> (others=>'0')));
    MULTS_5_37<=((others=> (others=>'0')));
    MULTS_5_38<=((others=> (others=>'0')));
    MULTS_5_39<=((others=> (others=>'0')));
    MULTS_5_40<=((others=> (others=>'0')));
    MULTS_5_41<=((others=> (others=>'0')));
    MULTS_5_42<=((others=> (others=>'0')));
    MULTS_5_43<=((others=> (others=>'0')));
    MULTS_5_44<=((others=> (others=>'0')));
    MULTS_5_45<=((others=> (others=>'0')));
    MULTS_5_46<=((others=> (others=>'0')));
    MULTS_5_47<=((others=> (others=>'0')));
    MULTS_5_48<=((others=> (others=>'0')));
    MULTS_5_49<=((others=> (others=>'0')));
    MULTS_5_50<=((others=> (others=>'0')));
    MULTS_5_51<=((others=> (others=>'0')));
    MULTS_5_52<=((others=> (others=>'0')));
    MULTS_5_53<=((others=> (others=>'0')));
    MULTS_5_54<=((others=> (others=>'0')));
    MULTS_5_55<=((others=> (others=>'0')));
    MULTS_5_56<=((others=> (others=>'0')));
    MULTS_5_57<=((others=> (others=>'0')));
    MULTS_5_58<=((others=> (others=>'0')));
    MULTS_5_59<=((others=> (others=>'0')));
    MULTS_5_60<=((others=> (others=>'0')));
    MULTS_5_61<=((others=> (others=>'0')));
    MULTS_5_62<=((others=> (others=>'0')));
    MULTS_5_63<=((others=> (others=>'0')));
    MULTS_5_64<=((others=> (others=>'0')));
    MULTS_5_65<=((others=> (others=>'0')));
    MULTS_5_66<=((others=> (others=>'0')));
    MULTS_5_67<=((others=> (others=>'0')));
    MULTS_5_68<=((others=> (others=>'0')));
    MULTS_5_69<=((others=> (others=>'0')));
    MULTS_5_70<=((others=> (others=>'0')));
    MULTS_5_71<=((others=> (others=>'0')));
    MULTS_5_72<=((others=> (others=>'0')));
    MULTS_5_73<=((others=> (others=>'0')));
    MULTS_5_74<=((others=> (others=>'0')));
    MULTS_5_75<=((others=> (others=>'0')));
    MULTS_5_76<=((others=> (others=>'0')));
    MULTS_5_77<=((others=> (others=>'0')));
    MULTS_5_78<=((others=> (others=>'0')));
    MULTS_5_79<=((others=> (others=>'0')));
    MULTS_5_80<=((others=> (others=>'0')));
    MULTS_5_81<=((others=> (others=>'0')));
    MULTS_5_82<=((others=> (others=>'0')));
    MULTS_5_83<=((others=> (others=>'0')));
    MULTS_5_84<=((others=> (others=>'0')));
    MULTS_5_85<=((others=> (others=>'0')));
    MULTS_5_86<=((others=> (others=>'0')));
    MULTS_5_87<=((others=> (others=>'0')));
    MULTS_5_88<=((others=> (others=>'0')));
    MULTS_5_89<=((others=> (others=>'0')));
    MULTS_5_90<=((others=> (others=>'0')));
    MULTS_5_91<=((others=> (others=>'0')));
    MULTS_5_92<=((others=> (others=>'0')));
    MULTS_5_93<=((others=> (others=>'0')));
    MULTS_5_94<=((others=> (others=>'0')));
    MULTS_5_95<=((others=> (others=>'0')));
    MULTS_5_96<=((others=> (others=>'0')));
    MULTS_5_97<=((others=> (others=>'0')));
    MULTS_5_98<=((others=> (others=>'0')));
    MULTS_5_99<=((others=> (others=>'0')));
    MULTS_5_100<=((others=> (others=>'0')));
    MULTS_5_101<=((others=> (others=>'0')));
    MULTS_5_102<=((others=> (others=>'0')));
    MULTS_5_103<=((others=> (others=>'0')));
    MULTS_5_104<=((others=> (others=>'0')));
    MULTS_5_105<=((others=> (others=>'0')));
    MULTS_5_106<=((others=> (others=>'0')));
    MULTS_5_107<=((others=> (others=>'0')));
    MULTS_5_108<=((others=> (others=>'0')));
    MULTS_5_109<=((others=> (others=>'0')));
    MULTS_5_110<=((others=> (others=>'0')));
    MULTS_5_111<=((others=> (others=>'0')));
    MULTS_5_112<=((others=> (others=>'0')));
    MULTS_5_113<=((others=> (others=>'0')));
    MULTS_5_114<=((others=> (others=>'0')));
    MULTS_5_115<=((others=> (others=>'0')));
    MULTS_5_116<=((others=> (others=>'0')));
    MULTS_5_117<=((others=> (others=>'0')));
    MULTS_5_118<=((others=> (others=>'0')));
    MULTS_5_119<=((others=> (others=>'0')));
    MULTS_5_120<=((others=> (others=>'0')));
    EN_SUM_MULT_6<='0';
    MULTS_6_1<=((others=> (others=>'0')));
    MULTS_6_2<=((others=> (others=>'0')));
    MULTS_6_3<=((others=> (others=>'0')));
    MULTS_6_4<=((others=> (others=>'0')));
    MULTS_6_5<=((others=> (others=>'0')));
    MULTS_6_6<=((others=> (others=>'0')));
    MULTS_6_7<=((others=> (others=>'0')));
    MULTS_6_8<=((others=> (others=>'0')));
    MULTS_6_9<=((others=> (others=>'0')));
    MULTS_6_10<=((others=> (others=>'0')));
    MULTS_6_11<=((others=> (others=>'0')));
    MULTS_6_12<=((others=> (others=>'0')));
    MULTS_6_13<=((others=> (others=>'0')));
    MULTS_6_14<=((others=> (others=>'0')));
    MULTS_6_15<=((others=> (others=>'0')));
    MULTS_6_16<=((others=> (others=>'0')));
    MULTS_6_17<=((others=> (others=>'0')));
    MULTS_6_18<=((others=> (others=>'0')));
    MULTS_6_19<=((others=> (others=>'0')));
    MULTS_6_20<=((others=> (others=>'0')));
    MULTS_6_21<=((others=> (others=>'0')));
    MULTS_6_22<=((others=> (others=>'0')));
    MULTS_6_23<=((others=> (others=>'0')));
    MULTS_6_24<=((others=> (others=>'0')));
    MULTS_6_25<=((others=> (others=>'0')));
    MULTS_6_26<=((others=> (others=>'0')));
    MULTS_6_27<=((others=> (others=>'0')));
    MULTS_6_28<=((others=> (others=>'0')));
    MULTS_6_29<=((others=> (others=>'0')));
    MULTS_6_30<=((others=> (others=>'0')));
    MULTS_6_31<=((others=> (others=>'0')));
    MULTS_6_32<=((others=> (others=>'0')));
    MULTS_6_33<=((others=> (others=>'0')));
    MULTS_6_34<=((others=> (others=>'0')));
    MULTS_6_35<=((others=> (others=>'0')));
    MULTS_6_36<=((others=> (others=>'0')));
    MULTS_6_37<=((others=> (others=>'0')));
    MULTS_6_38<=((others=> (others=>'0')));
    MULTS_6_39<=((others=> (others=>'0')));
    MULTS_6_40<=((others=> (others=>'0')));
    MULTS_6_41<=((others=> (others=>'0')));
    MULTS_6_42<=((others=> (others=>'0')));
    MULTS_6_43<=((others=> (others=>'0')));
    MULTS_6_44<=((others=> (others=>'0')));
    MULTS_6_45<=((others=> (others=>'0')));
    MULTS_6_46<=((others=> (others=>'0')));
    MULTS_6_47<=((others=> (others=>'0')));
    MULTS_6_48<=((others=> (others=>'0')));
    MULTS_6_49<=((others=> (others=>'0')));
    MULTS_6_50<=((others=> (others=>'0')));
    MULTS_6_51<=((others=> (others=>'0')));
    MULTS_6_52<=((others=> (others=>'0')));
    MULTS_6_53<=((others=> (others=>'0')));
    MULTS_6_54<=((others=> (others=>'0')));
    MULTS_6_55<=((others=> (others=>'0')));
    MULTS_6_56<=((others=> (others=>'0')));
    MULTS_6_57<=((others=> (others=>'0')));
    MULTS_6_58<=((others=> (others=>'0')));
    MULTS_6_59<=((others=> (others=>'0')));
    MULTS_6_60<=((others=> (others=>'0')));
    MULTS_6_61<=((others=> (others=>'0')));
    MULTS_6_62<=((others=> (others=>'0')));
    MULTS_6_63<=((others=> (others=>'0')));
    MULTS_6_64<=((others=> (others=>'0')));
    MULTS_6_65<=((others=> (others=>'0')));
    MULTS_6_66<=((others=> (others=>'0')));
    MULTS_6_67<=((others=> (others=>'0')));
    MULTS_6_68<=((others=> (others=>'0')));
    MULTS_6_69<=((others=> (others=>'0')));
    MULTS_6_70<=((others=> (others=>'0')));
    MULTS_6_71<=((others=> (others=>'0')));
    MULTS_6_72<=((others=> (others=>'0')));
    MULTS_6_73<=((others=> (others=>'0')));
    MULTS_6_74<=((others=> (others=>'0')));
    MULTS_6_75<=((others=> (others=>'0')));
    MULTS_6_76<=((others=> (others=>'0')));
    MULTS_6_77<=((others=> (others=>'0')));
    MULTS_6_78<=((others=> (others=>'0')));
    MULTS_6_79<=((others=> (others=>'0')));
    MULTS_6_80<=((others=> (others=>'0')));
    MULTS_6_81<=((others=> (others=>'0')));
    MULTS_6_82<=((others=> (others=>'0')));
    MULTS_6_83<=((others=> (others=>'0')));
    MULTS_6_84<=((others=> (others=>'0')));
    MULTS_6_85<=((others=> (others=>'0')));
    MULTS_6_86<=((others=> (others=>'0')));
    MULTS_6_87<=((others=> (others=>'0')));
    MULTS_6_88<=((others=> (others=>'0')));
    MULTS_6_89<=((others=> (others=>'0')));
    MULTS_6_90<=((others=> (others=>'0')));
    MULTS_6_91<=((others=> (others=>'0')));
    MULTS_6_92<=((others=> (others=>'0')));
    MULTS_6_93<=((others=> (others=>'0')));
    MULTS_6_94<=((others=> (others=>'0')));
    MULTS_6_95<=((others=> (others=>'0')));
    MULTS_6_96<=((others=> (others=>'0')));
    MULTS_6_97<=((others=> (others=>'0')));
    MULTS_6_98<=((others=> (others=>'0')));
    MULTS_6_99<=((others=> (others=>'0')));
    MULTS_6_100<=((others=> (others=>'0')));
    MULTS_6_101<=((others=> (others=>'0')));
    MULTS_6_102<=((others=> (others=>'0')));
    MULTS_6_103<=((others=> (others=>'0')));
    MULTS_6_104<=((others=> (others=>'0')));
    MULTS_6_105<=((others=> (others=>'0')));
    MULTS_6_106<=((others=> (others=>'0')));
    MULTS_6_107<=((others=> (others=>'0')));
    MULTS_6_108<=((others=> (others=>'0')));
    MULTS_6_109<=((others=> (others=>'0')));
    MULTS_6_110<=((others=> (others=>'0')));
    MULTS_6_111<=((others=> (others=>'0')));
    MULTS_6_112<=((others=> (others=>'0')));
    MULTS_6_113<=((others=> (others=>'0')));
    MULTS_6_114<=((others=> (others=>'0')));
    MULTS_6_115<=((others=> (others=>'0')));
    MULTS_6_116<=((others=> (others=>'0')));
    MULTS_6_117<=((others=> (others=>'0')));
    MULTS_6_118<=((others=> (others=>'0')));
    MULTS_6_119<=((others=> (others=>'0')));
    MULTS_6_120<=((others=> (others=>'0')));
    EN_SUM_MULT_7<='0';
    MULTS_7_1<=((others=> (others=>'0')));
    MULTS_7_2<=((others=> (others=>'0')));
    MULTS_7_3<=((others=> (others=>'0')));
    MULTS_7_4<=((others=> (others=>'0')));
    MULTS_7_5<=((others=> (others=>'0')));
    MULTS_7_6<=((others=> (others=>'0')));
    MULTS_7_7<=((others=> (others=>'0')));
    MULTS_7_8<=((others=> (others=>'0')));
    MULTS_7_9<=((others=> (others=>'0')));
    MULTS_7_10<=((others=> (others=>'0')));
    MULTS_7_11<=((others=> (others=>'0')));
    MULTS_7_12<=((others=> (others=>'0')));
    MULTS_7_13<=((others=> (others=>'0')));
    MULTS_7_14<=((others=> (others=>'0')));
    MULTS_7_15<=((others=> (others=>'0')));
    MULTS_7_16<=((others=> (others=>'0')));
    MULTS_7_17<=((others=> (others=>'0')));
    MULTS_7_18<=((others=> (others=>'0')));
    MULTS_7_19<=((others=> (others=>'0')));
    MULTS_7_20<=((others=> (others=>'0')));
    MULTS_7_21<=((others=> (others=>'0')));
    MULTS_7_22<=((others=> (others=>'0')));
    MULTS_7_23<=((others=> (others=>'0')));
    MULTS_7_24<=((others=> (others=>'0')));
    MULTS_7_25<=((others=> (others=>'0')));
    MULTS_7_26<=((others=> (others=>'0')));
    MULTS_7_27<=((others=> (others=>'0')));
    MULTS_7_28<=((others=> (others=>'0')));
    MULTS_7_29<=((others=> (others=>'0')));
    MULTS_7_30<=((others=> (others=>'0')));
    MULTS_7_31<=((others=> (others=>'0')));
    MULTS_7_32<=((others=> (others=>'0')));
    MULTS_7_33<=((others=> (others=>'0')));
    MULTS_7_34<=((others=> (others=>'0')));
    MULTS_7_35<=((others=> (others=>'0')));
    MULTS_7_36<=((others=> (others=>'0')));
    MULTS_7_37<=((others=> (others=>'0')));
    MULTS_7_38<=((others=> (others=>'0')));
    MULTS_7_39<=((others=> (others=>'0')));
    MULTS_7_40<=((others=> (others=>'0')));
    MULTS_7_41<=((others=> (others=>'0')));
    MULTS_7_42<=((others=> (others=>'0')));
    MULTS_7_43<=((others=> (others=>'0')));
    MULTS_7_44<=((others=> (others=>'0')));
    MULTS_7_45<=((others=> (others=>'0')));
    MULTS_7_46<=((others=> (others=>'0')));
    MULTS_7_47<=((others=> (others=>'0')));
    MULTS_7_48<=((others=> (others=>'0')));
    MULTS_7_49<=((others=> (others=>'0')));
    MULTS_7_50<=((others=> (others=>'0')));
    MULTS_7_51<=((others=> (others=>'0')));
    MULTS_7_52<=((others=> (others=>'0')));
    MULTS_7_53<=((others=> (others=>'0')));
    MULTS_7_54<=((others=> (others=>'0')));
    MULTS_7_55<=((others=> (others=>'0')));
    MULTS_7_56<=((others=> (others=>'0')));
    MULTS_7_57<=((others=> (others=>'0')));
    MULTS_7_58<=((others=> (others=>'0')));
    MULTS_7_59<=((others=> (others=>'0')));
    MULTS_7_60<=((others=> (others=>'0')));
    MULTS_7_61<=((others=> (others=>'0')));
    MULTS_7_62<=((others=> (others=>'0')));
    MULTS_7_63<=((others=> (others=>'0')));
    MULTS_7_64<=((others=> (others=>'0')));
    MULTS_7_65<=((others=> (others=>'0')));
    MULTS_7_66<=((others=> (others=>'0')));
    MULTS_7_67<=((others=> (others=>'0')));
    MULTS_7_68<=((others=> (others=>'0')));
    MULTS_7_69<=((others=> (others=>'0')));
    MULTS_7_70<=((others=> (others=>'0')));
    MULTS_7_71<=((others=> (others=>'0')));
    MULTS_7_72<=((others=> (others=>'0')));
    MULTS_7_73<=((others=> (others=>'0')));
    MULTS_7_74<=((others=> (others=>'0')));
    MULTS_7_75<=((others=> (others=>'0')));
    MULTS_7_76<=((others=> (others=>'0')));
    MULTS_7_77<=((others=> (others=>'0')));
    MULTS_7_78<=((others=> (others=>'0')));
    MULTS_7_79<=((others=> (others=>'0')));
    MULTS_7_80<=((others=> (others=>'0')));
    MULTS_7_81<=((others=> (others=>'0')));
    MULTS_7_82<=((others=> (others=>'0')));
    MULTS_7_83<=((others=> (others=>'0')));
    MULTS_7_84<=((others=> (others=>'0')));
    MULTS_7_85<=((others=> (others=>'0')));
    MULTS_7_86<=((others=> (others=>'0')));
    MULTS_7_87<=((others=> (others=>'0')));
    MULTS_7_88<=((others=> (others=>'0')));
    MULTS_7_89<=((others=> (others=>'0')));
    MULTS_7_90<=((others=> (others=>'0')));
    MULTS_7_91<=((others=> (others=>'0')));
    MULTS_7_92<=((others=> (others=>'0')));
    MULTS_7_93<=((others=> (others=>'0')));
    MULTS_7_94<=((others=> (others=>'0')));
    MULTS_7_95<=((others=> (others=>'0')));
    MULTS_7_96<=((others=> (others=>'0')));
    MULTS_7_97<=((others=> (others=>'0')));
    MULTS_7_98<=((others=> (others=>'0')));
    MULTS_7_99<=((others=> (others=>'0')));
    MULTS_7_100<=((others=> (others=>'0')));
    MULTS_7_101<=((others=> (others=>'0')));
    MULTS_7_102<=((others=> (others=>'0')));
    MULTS_7_103<=((others=> (others=>'0')));
    MULTS_7_104<=((others=> (others=>'0')));
    MULTS_7_105<=((others=> (others=>'0')));
    MULTS_7_106<=((others=> (others=>'0')));
    MULTS_7_107<=((others=> (others=>'0')));
    MULTS_7_108<=((others=> (others=>'0')));
    MULTS_7_109<=((others=> (others=>'0')));
    MULTS_7_110<=((others=> (others=>'0')));
    MULTS_7_111<=((others=> (others=>'0')));
    MULTS_7_112<=((others=> (others=>'0')));
    MULTS_7_113<=((others=> (others=>'0')));
    MULTS_7_114<=((others=> (others=>'0')));
    MULTS_7_115<=((others=> (others=>'0')));
    MULTS_7_116<=((others=> (others=>'0')));
    MULTS_7_117<=((others=> (others=>'0')));
    MULTS_7_118<=((others=> (others=>'0')));
    MULTS_7_119<=((others=> (others=>'0')));
    MULTS_7_120<=((others=> (others=>'0')));

------------------------------------------------ PROCESS START------------------------------------------------------
	  
   else 	
	if EN_LOC_STREAM_7='1' and EN_STREAM= '1' and OUT_PIXEL_COUNT<VALID_CYCLES  then    -- check valid data and enable stream
		
		if  FRST_TIM_EN_7='1' then EN_NXT_LYR_7<='1';end if;

			MULT_1(0)<=signed(DIN_1_7)*signed(FMAP_1_1);
			MULT_2(0)<=signed(DIN_2_7)*signed(FMAP_1_2);
			MULT_3(0)<=signed(DIN_3_7)*signed(FMAP_1_3);
			MULT_4(0)<=signed(DIN_4_7)*signed(FMAP_1_4);
			MULT_5(0)<=signed(DIN_5_7)*signed(FMAP_1_5);
			MULT_6(0)<=signed(DIN_6_7)*signed(FMAP_1_6);
			MULT_7(0)<=signed(DIN_7_7)*signed(FMAP_1_7);
			MULT_8(0)<=signed(DIN_8_7)*signed(FMAP_1_8);
			MULT_9(0)<=signed(DIN_9_7)*signed(FMAP_1_9);
			MULT_10(0)<=signed(DIN_10_7)*signed(FMAP_1_10);
			MULT_11(0)<=signed(DIN_11_7)*signed(FMAP_1_11);
			MULT_12(0)<=signed(DIN_12_7)*signed(FMAP_1_12);
			MULT_13(0)<=signed(DIN_13_7)*signed(FMAP_1_13);
			MULT_14(0)<=signed(DIN_14_7)*signed(FMAP_1_14);
			MULT_15(0)<=signed(DIN_15_7)*signed(FMAP_1_15);
			MULT_16(0)<=signed(DIN_16_7)*signed(FMAP_1_16);
			MULT_17(0)<=signed(DIN_17_7)*signed(FMAP_1_17);
			MULT_18(0)<=signed(DIN_18_7)*signed(FMAP_1_18);
			MULT_19(0)<=signed(DIN_19_7)*signed(FMAP_1_19);
			MULT_20(0)<=signed(DIN_20_7)*signed(FMAP_1_20);
			MULT_21(0)<=signed(DIN_21_7)*signed(FMAP_1_21);
			MULT_22(0)<=signed(DIN_22_7)*signed(FMAP_1_22);
			MULT_23(0)<=signed(DIN_23_7)*signed(FMAP_1_23);
			MULT_24(0)<=signed(DIN_24_7)*signed(FMAP_1_24);
			MULT_25(0)<=signed(DIN_25_7)*signed(FMAP_1_25);
			MULT_26(0)<=signed(DIN_26_7)*signed(FMAP_1_26);
			MULT_27(0)<=signed(DIN_27_7)*signed(FMAP_1_27);
			MULT_28(0)<=signed(DIN_28_7)*signed(FMAP_1_28);
			MULT_29(0)<=signed(DIN_29_7)*signed(FMAP_1_29);
			MULT_30(0)<=signed(DIN_30_7)*signed(FMAP_1_30);
			MULT_31(0)<=signed(DIN_31_7)*signed(FMAP_1_31);
			MULT_32(0)<=signed(DIN_32_7)*signed(FMAP_1_32);
			MULT_33(0)<=signed(DIN_33_7)*signed(FMAP_1_33);
			MULT_34(0)<=signed(DIN_34_7)*signed(FMAP_1_34);
			MULT_35(0)<=signed(DIN_35_7)*signed(FMAP_1_35);
			MULT_36(0)<=signed(DIN_36_7)*signed(FMAP_1_36);
			MULT_37(0)<=signed(DIN_37_7)*signed(FMAP_1_37);
			MULT_38(0)<=signed(DIN_38_7)*signed(FMAP_1_38);
			MULT_39(0)<=signed(DIN_39_7)*signed(FMAP_1_39);
			MULT_40(0)<=signed(DIN_40_7)*signed(FMAP_1_40);
			MULT_41(0)<=signed(DIN_41_7)*signed(FMAP_1_41);
			MULT_42(0)<=signed(DIN_42_7)*signed(FMAP_1_42);
			MULT_43(0)<=signed(DIN_43_7)*signed(FMAP_1_43);
			MULT_44(0)<=signed(DIN_44_7)*signed(FMAP_1_44);
			MULT_45(0)<=signed(DIN_45_7)*signed(FMAP_1_45);
			MULT_46(0)<=signed(DIN_46_7)*signed(FMAP_1_46);
			MULT_47(0)<=signed(DIN_47_7)*signed(FMAP_1_47);
			MULT_48(0)<=signed(DIN_48_7)*signed(FMAP_1_48);
			MULT_49(0)<=signed(DIN_49_7)*signed(FMAP_1_49);
			MULT_50(0)<=signed(DIN_50_7)*signed(FMAP_1_50);
			MULT_51(0)<=signed(DIN_51_7)*signed(FMAP_1_51);
			MULT_52(0)<=signed(DIN_52_7)*signed(FMAP_1_52);
			MULT_53(0)<=signed(DIN_53_7)*signed(FMAP_1_53);
			MULT_54(0)<=signed(DIN_54_7)*signed(FMAP_1_54);
			MULT_55(0)<=signed(DIN_55_7)*signed(FMAP_1_55);
			MULT_56(0)<=signed(DIN_56_7)*signed(FMAP_1_56);
			MULT_57(0)<=signed(DIN_57_7)*signed(FMAP_1_57);
			MULT_58(0)<=signed(DIN_58_7)*signed(FMAP_1_58);
			MULT_59(0)<=signed(DIN_59_7)*signed(FMAP_1_59);
			MULT_60(0)<=signed(DIN_60_7)*signed(FMAP_1_60);
			MULT_61(0)<=signed(DIN_61_7)*signed(FMAP_1_61);
			MULT_62(0)<=signed(DIN_62_7)*signed(FMAP_1_62);
			MULT_63(0)<=signed(DIN_63_7)*signed(FMAP_1_63);
			MULT_64(0)<=signed(DIN_64_7)*signed(FMAP_1_64);
			MULT_65(0)<=signed(DIN_65_7)*signed(FMAP_1_65);
			MULT_66(0)<=signed(DIN_66_7)*signed(FMAP_1_66);
			MULT_67(0)<=signed(DIN_67_7)*signed(FMAP_1_67);
			MULT_68(0)<=signed(DIN_68_7)*signed(FMAP_1_68);
			MULT_69(0)<=signed(DIN_69_7)*signed(FMAP_1_69);
			MULT_70(0)<=signed(DIN_70_7)*signed(FMAP_1_70);
			MULT_71(0)<=signed(DIN_71_7)*signed(FMAP_1_71);
			MULT_72(0)<=signed(DIN_72_7)*signed(FMAP_1_72);
			MULT_73(0)<=signed(DIN_73_7)*signed(FMAP_1_73);
			MULT_74(0)<=signed(DIN_74_7)*signed(FMAP_1_74);
			MULT_75(0)<=signed(DIN_75_7)*signed(FMAP_1_75);
			MULT_76(0)<=signed(DIN_76_7)*signed(FMAP_1_76);
			MULT_77(0)<=signed(DIN_77_7)*signed(FMAP_1_77);
			MULT_78(0)<=signed(DIN_78_7)*signed(FMAP_1_78);
			MULT_79(0)<=signed(DIN_79_7)*signed(FMAP_1_79);
			MULT_80(0)<=signed(DIN_80_7)*signed(FMAP_1_80);
			MULT_81(0)<=signed(DIN_81_7)*signed(FMAP_1_81);
			MULT_82(0)<=signed(DIN_82_7)*signed(FMAP_1_82);
			MULT_83(0)<=signed(DIN_83_7)*signed(FMAP_1_83);
			MULT_84(0)<=signed(DIN_84_7)*signed(FMAP_1_84);
			MULT_85(0)<=signed(DIN_85_7)*signed(FMAP_1_85);
			MULT_86(0)<=signed(DIN_86_7)*signed(FMAP_1_86);
			MULT_87(0)<=signed(DIN_87_7)*signed(FMAP_1_87);
			MULT_88(0)<=signed(DIN_88_7)*signed(FMAP_1_88);
			MULT_89(0)<=signed(DIN_89_7)*signed(FMAP_1_89);
			MULT_90(0)<=signed(DIN_90_7)*signed(FMAP_1_90);
			MULT_91(0)<=signed(DIN_91_7)*signed(FMAP_1_91);
			MULT_92(0)<=signed(DIN_92_7)*signed(FMAP_1_92);
			MULT_93(0)<=signed(DIN_93_7)*signed(FMAP_1_93);
			MULT_94(0)<=signed(DIN_94_7)*signed(FMAP_1_94);
			MULT_95(0)<=signed(DIN_95_7)*signed(FMAP_1_95);
			MULT_96(0)<=signed(DIN_96_7)*signed(FMAP_1_96);
			MULT_97(0)<=signed(DIN_97_7)*signed(FMAP_1_97);
			MULT_98(0)<=signed(DIN_98_7)*signed(FMAP_1_98);
			MULT_99(0)<=signed(DIN_99_7)*signed(FMAP_1_99);
			MULT_100(0)<=signed(DIN_100_7)*signed(FMAP_1_100);
			MULT_101(0)<=signed(DIN_101_7)*signed(FMAP_1_101);
			MULT_102(0)<=signed(DIN_102_7)*signed(FMAP_1_102);
			MULT_103(0)<=signed(DIN_103_7)*signed(FMAP_1_103);
			MULT_104(0)<=signed(DIN_104_7)*signed(FMAP_1_104);
			MULT_105(0)<=signed(DIN_105_7)*signed(FMAP_1_105);
			MULT_106(0)<=signed(DIN_106_7)*signed(FMAP_1_106);
			MULT_107(0)<=signed(DIN_107_7)*signed(FMAP_1_107);
			MULT_108(0)<=signed(DIN_108_7)*signed(FMAP_1_108);
			MULT_109(0)<=signed(DIN_109_7)*signed(FMAP_1_109);
			MULT_110(0)<=signed(DIN_110_7)*signed(FMAP_1_110);
			MULT_111(0)<=signed(DIN_111_7)*signed(FMAP_1_111);
			MULT_112(0)<=signed(DIN_112_7)*signed(FMAP_1_112);
			MULT_113(0)<=signed(DIN_113_7)*signed(FMAP_1_113);
			MULT_114(0)<=signed(DIN_114_7)*signed(FMAP_1_114);
			MULT_115(0)<=signed(DIN_115_7)*signed(FMAP_1_115);
			MULT_116(0)<=signed(DIN_116_7)*signed(FMAP_1_116);
			MULT_117(0)<=signed(DIN_117_7)*signed(FMAP_1_117);
			MULT_118(0)<=signed(DIN_118_7)*signed(FMAP_1_118);
			MULT_119(0)<=signed(DIN_119_7)*signed(FMAP_1_119);
			MULT_120(0)<=signed(DIN_120_7)*signed(FMAP_1_120);

			MULT_1(1)<=signed(DIN_1_7)*signed(FMAP_2_1);
			MULT_2(1)<=signed(DIN_2_7)*signed(FMAP_2_2);
			MULT_3(1)<=signed(DIN_3_7)*signed(FMAP_2_3);
			MULT_4(1)<=signed(DIN_4_7)*signed(FMAP_2_4);
			MULT_5(1)<=signed(DIN_5_7)*signed(FMAP_2_5);
			MULT_6(1)<=signed(DIN_6_7)*signed(FMAP_2_6);
			MULT_7(1)<=signed(DIN_7_7)*signed(FMAP_2_7);
			MULT_8(1)<=signed(DIN_8_7)*signed(FMAP_2_8);
			MULT_9(1)<=signed(DIN_9_7)*signed(FMAP_2_9);
			MULT_10(1)<=signed(DIN_10_7)*signed(FMAP_2_10);
			MULT_11(1)<=signed(DIN_11_7)*signed(FMAP_2_11);
			MULT_12(1)<=signed(DIN_12_7)*signed(FMAP_2_12);
			MULT_13(1)<=signed(DIN_13_7)*signed(FMAP_2_13);
			MULT_14(1)<=signed(DIN_14_7)*signed(FMAP_2_14);
			MULT_15(1)<=signed(DIN_15_7)*signed(FMAP_2_15);
			MULT_16(1)<=signed(DIN_16_7)*signed(FMAP_2_16);
			MULT_17(1)<=signed(DIN_17_7)*signed(FMAP_2_17);
			MULT_18(1)<=signed(DIN_18_7)*signed(FMAP_2_18);
			MULT_19(1)<=signed(DIN_19_7)*signed(FMAP_2_19);
			MULT_20(1)<=signed(DIN_20_7)*signed(FMAP_2_20);
			MULT_21(1)<=signed(DIN_21_7)*signed(FMAP_2_21);
			MULT_22(1)<=signed(DIN_22_7)*signed(FMAP_2_22);
			MULT_23(1)<=signed(DIN_23_7)*signed(FMAP_2_23);
			MULT_24(1)<=signed(DIN_24_7)*signed(FMAP_2_24);
			MULT_25(1)<=signed(DIN_25_7)*signed(FMAP_2_25);
			MULT_26(1)<=signed(DIN_26_7)*signed(FMAP_2_26);
			MULT_27(1)<=signed(DIN_27_7)*signed(FMAP_2_27);
			MULT_28(1)<=signed(DIN_28_7)*signed(FMAP_2_28);
			MULT_29(1)<=signed(DIN_29_7)*signed(FMAP_2_29);
			MULT_30(1)<=signed(DIN_30_7)*signed(FMAP_2_30);
			MULT_31(1)<=signed(DIN_31_7)*signed(FMAP_2_31);
			MULT_32(1)<=signed(DIN_32_7)*signed(FMAP_2_32);
			MULT_33(1)<=signed(DIN_33_7)*signed(FMAP_2_33);
			MULT_34(1)<=signed(DIN_34_7)*signed(FMAP_2_34);
			MULT_35(1)<=signed(DIN_35_7)*signed(FMAP_2_35);
			MULT_36(1)<=signed(DIN_36_7)*signed(FMAP_2_36);
			MULT_37(1)<=signed(DIN_37_7)*signed(FMAP_2_37);
			MULT_38(1)<=signed(DIN_38_7)*signed(FMAP_2_38);
			MULT_39(1)<=signed(DIN_39_7)*signed(FMAP_2_39);
			MULT_40(1)<=signed(DIN_40_7)*signed(FMAP_2_40);
			MULT_41(1)<=signed(DIN_41_7)*signed(FMAP_2_41);
			MULT_42(1)<=signed(DIN_42_7)*signed(FMAP_2_42);
			MULT_43(1)<=signed(DIN_43_7)*signed(FMAP_2_43);
			MULT_44(1)<=signed(DIN_44_7)*signed(FMAP_2_44);
			MULT_45(1)<=signed(DIN_45_7)*signed(FMAP_2_45);
			MULT_46(1)<=signed(DIN_46_7)*signed(FMAP_2_46);
			MULT_47(1)<=signed(DIN_47_7)*signed(FMAP_2_47);
			MULT_48(1)<=signed(DIN_48_7)*signed(FMAP_2_48);
			MULT_49(1)<=signed(DIN_49_7)*signed(FMAP_2_49);
			MULT_50(1)<=signed(DIN_50_7)*signed(FMAP_2_50);
			MULT_51(1)<=signed(DIN_51_7)*signed(FMAP_2_51);
			MULT_52(1)<=signed(DIN_52_7)*signed(FMAP_2_52);
			MULT_53(1)<=signed(DIN_53_7)*signed(FMAP_2_53);
			MULT_54(1)<=signed(DIN_54_7)*signed(FMAP_2_54);
			MULT_55(1)<=signed(DIN_55_7)*signed(FMAP_2_55);
			MULT_56(1)<=signed(DIN_56_7)*signed(FMAP_2_56);
			MULT_57(1)<=signed(DIN_57_7)*signed(FMAP_2_57);
			MULT_58(1)<=signed(DIN_58_7)*signed(FMAP_2_58);
			MULT_59(1)<=signed(DIN_59_7)*signed(FMAP_2_59);
			MULT_60(1)<=signed(DIN_60_7)*signed(FMAP_2_60);
			MULT_61(1)<=signed(DIN_61_7)*signed(FMAP_2_61);
			MULT_62(1)<=signed(DIN_62_7)*signed(FMAP_2_62);
			MULT_63(1)<=signed(DIN_63_7)*signed(FMAP_2_63);
			MULT_64(1)<=signed(DIN_64_7)*signed(FMAP_2_64);
			MULT_65(1)<=signed(DIN_65_7)*signed(FMAP_2_65);
			MULT_66(1)<=signed(DIN_66_7)*signed(FMAP_2_66);
			MULT_67(1)<=signed(DIN_67_7)*signed(FMAP_2_67);
			MULT_68(1)<=signed(DIN_68_7)*signed(FMAP_2_68);
			MULT_69(1)<=signed(DIN_69_7)*signed(FMAP_2_69);
			MULT_70(1)<=signed(DIN_70_7)*signed(FMAP_2_70);
			MULT_71(1)<=signed(DIN_71_7)*signed(FMAP_2_71);
			MULT_72(1)<=signed(DIN_72_7)*signed(FMAP_2_72);
			MULT_73(1)<=signed(DIN_73_7)*signed(FMAP_2_73);
			MULT_74(1)<=signed(DIN_74_7)*signed(FMAP_2_74);
			MULT_75(1)<=signed(DIN_75_7)*signed(FMAP_2_75);
			MULT_76(1)<=signed(DIN_76_7)*signed(FMAP_2_76);
			MULT_77(1)<=signed(DIN_77_7)*signed(FMAP_2_77);
			MULT_78(1)<=signed(DIN_78_7)*signed(FMAP_2_78);
			MULT_79(1)<=signed(DIN_79_7)*signed(FMAP_2_79);
			MULT_80(1)<=signed(DIN_80_7)*signed(FMAP_2_80);
			MULT_81(1)<=signed(DIN_81_7)*signed(FMAP_2_81);
			MULT_82(1)<=signed(DIN_82_7)*signed(FMAP_2_82);
			MULT_83(1)<=signed(DIN_83_7)*signed(FMAP_2_83);
			MULT_84(1)<=signed(DIN_84_7)*signed(FMAP_2_84);
			MULT_85(1)<=signed(DIN_85_7)*signed(FMAP_2_85);
			MULT_86(1)<=signed(DIN_86_7)*signed(FMAP_2_86);
			MULT_87(1)<=signed(DIN_87_7)*signed(FMAP_2_87);
			MULT_88(1)<=signed(DIN_88_7)*signed(FMAP_2_88);
			MULT_89(1)<=signed(DIN_89_7)*signed(FMAP_2_89);
			MULT_90(1)<=signed(DIN_90_7)*signed(FMAP_2_90);
			MULT_91(1)<=signed(DIN_91_7)*signed(FMAP_2_91);
			MULT_92(1)<=signed(DIN_92_7)*signed(FMAP_2_92);
			MULT_93(1)<=signed(DIN_93_7)*signed(FMAP_2_93);
			MULT_94(1)<=signed(DIN_94_7)*signed(FMAP_2_94);
			MULT_95(1)<=signed(DIN_95_7)*signed(FMAP_2_95);
			MULT_96(1)<=signed(DIN_96_7)*signed(FMAP_2_96);
			MULT_97(1)<=signed(DIN_97_7)*signed(FMAP_2_97);
			MULT_98(1)<=signed(DIN_98_7)*signed(FMAP_2_98);
			MULT_99(1)<=signed(DIN_99_7)*signed(FMAP_2_99);
			MULT_100(1)<=signed(DIN_100_7)*signed(FMAP_2_100);
			MULT_101(1)<=signed(DIN_101_7)*signed(FMAP_2_101);
			MULT_102(1)<=signed(DIN_102_7)*signed(FMAP_2_102);
			MULT_103(1)<=signed(DIN_103_7)*signed(FMAP_2_103);
			MULT_104(1)<=signed(DIN_104_7)*signed(FMAP_2_104);
			MULT_105(1)<=signed(DIN_105_7)*signed(FMAP_2_105);
			MULT_106(1)<=signed(DIN_106_7)*signed(FMAP_2_106);
			MULT_107(1)<=signed(DIN_107_7)*signed(FMAP_2_107);
			MULT_108(1)<=signed(DIN_108_7)*signed(FMAP_2_108);
			MULT_109(1)<=signed(DIN_109_7)*signed(FMAP_2_109);
			MULT_110(1)<=signed(DIN_110_7)*signed(FMAP_2_110);
			MULT_111(1)<=signed(DIN_111_7)*signed(FMAP_2_111);
			MULT_112(1)<=signed(DIN_112_7)*signed(FMAP_2_112);
			MULT_113(1)<=signed(DIN_113_7)*signed(FMAP_2_113);
			MULT_114(1)<=signed(DIN_114_7)*signed(FMAP_2_114);
			MULT_115(1)<=signed(DIN_115_7)*signed(FMAP_2_115);
			MULT_116(1)<=signed(DIN_116_7)*signed(FMAP_2_116);
			MULT_117(1)<=signed(DIN_117_7)*signed(FMAP_2_117);
			MULT_118(1)<=signed(DIN_118_7)*signed(FMAP_2_118);
			MULT_119(1)<=signed(DIN_119_7)*signed(FMAP_2_119);
			MULT_120(1)<=signed(DIN_120_7)*signed(FMAP_2_120);

			MULT_1(2)<=signed(DIN_1_7)*signed(FMAP_3_1);
			MULT_2(2)<=signed(DIN_2_7)*signed(FMAP_3_2);
			MULT_3(2)<=signed(DIN_3_7)*signed(FMAP_3_3);
			MULT_4(2)<=signed(DIN_4_7)*signed(FMAP_3_4);
			MULT_5(2)<=signed(DIN_5_7)*signed(FMAP_3_5);
			MULT_6(2)<=signed(DIN_6_7)*signed(FMAP_3_6);
			MULT_7(2)<=signed(DIN_7_7)*signed(FMAP_3_7);
			MULT_8(2)<=signed(DIN_8_7)*signed(FMAP_3_8);
			MULT_9(2)<=signed(DIN_9_7)*signed(FMAP_3_9);
			MULT_10(2)<=signed(DIN_10_7)*signed(FMAP_3_10);
			MULT_11(2)<=signed(DIN_11_7)*signed(FMAP_3_11);
			MULT_12(2)<=signed(DIN_12_7)*signed(FMAP_3_12);
			MULT_13(2)<=signed(DIN_13_7)*signed(FMAP_3_13);
			MULT_14(2)<=signed(DIN_14_7)*signed(FMAP_3_14);
			MULT_15(2)<=signed(DIN_15_7)*signed(FMAP_3_15);
			MULT_16(2)<=signed(DIN_16_7)*signed(FMAP_3_16);
			MULT_17(2)<=signed(DIN_17_7)*signed(FMAP_3_17);
			MULT_18(2)<=signed(DIN_18_7)*signed(FMAP_3_18);
			MULT_19(2)<=signed(DIN_19_7)*signed(FMAP_3_19);
			MULT_20(2)<=signed(DIN_20_7)*signed(FMAP_3_20);
			MULT_21(2)<=signed(DIN_21_7)*signed(FMAP_3_21);
			MULT_22(2)<=signed(DIN_22_7)*signed(FMAP_3_22);
			MULT_23(2)<=signed(DIN_23_7)*signed(FMAP_3_23);
			MULT_24(2)<=signed(DIN_24_7)*signed(FMAP_3_24);
			MULT_25(2)<=signed(DIN_25_7)*signed(FMAP_3_25);
			MULT_26(2)<=signed(DIN_26_7)*signed(FMAP_3_26);
			MULT_27(2)<=signed(DIN_27_7)*signed(FMAP_3_27);
			MULT_28(2)<=signed(DIN_28_7)*signed(FMAP_3_28);
			MULT_29(2)<=signed(DIN_29_7)*signed(FMAP_3_29);
			MULT_30(2)<=signed(DIN_30_7)*signed(FMAP_3_30);
			MULT_31(2)<=signed(DIN_31_7)*signed(FMAP_3_31);
			MULT_32(2)<=signed(DIN_32_7)*signed(FMAP_3_32);
			MULT_33(2)<=signed(DIN_33_7)*signed(FMAP_3_33);
			MULT_34(2)<=signed(DIN_34_7)*signed(FMAP_3_34);
			MULT_35(2)<=signed(DIN_35_7)*signed(FMAP_3_35);
			MULT_36(2)<=signed(DIN_36_7)*signed(FMAP_3_36);
			MULT_37(2)<=signed(DIN_37_7)*signed(FMAP_3_37);
			MULT_38(2)<=signed(DIN_38_7)*signed(FMAP_3_38);
			MULT_39(2)<=signed(DIN_39_7)*signed(FMAP_3_39);
			MULT_40(2)<=signed(DIN_40_7)*signed(FMAP_3_40);
			MULT_41(2)<=signed(DIN_41_7)*signed(FMAP_3_41);
			MULT_42(2)<=signed(DIN_42_7)*signed(FMAP_3_42);
			MULT_43(2)<=signed(DIN_43_7)*signed(FMAP_3_43);
			MULT_44(2)<=signed(DIN_44_7)*signed(FMAP_3_44);
			MULT_45(2)<=signed(DIN_45_7)*signed(FMAP_3_45);
			MULT_46(2)<=signed(DIN_46_7)*signed(FMAP_3_46);
			MULT_47(2)<=signed(DIN_47_7)*signed(FMAP_3_47);
			MULT_48(2)<=signed(DIN_48_7)*signed(FMAP_3_48);
			MULT_49(2)<=signed(DIN_49_7)*signed(FMAP_3_49);
			MULT_50(2)<=signed(DIN_50_7)*signed(FMAP_3_50);
			MULT_51(2)<=signed(DIN_51_7)*signed(FMAP_3_51);
			MULT_52(2)<=signed(DIN_52_7)*signed(FMAP_3_52);
			MULT_53(2)<=signed(DIN_53_7)*signed(FMAP_3_53);
			MULT_54(2)<=signed(DIN_54_7)*signed(FMAP_3_54);
			MULT_55(2)<=signed(DIN_55_7)*signed(FMAP_3_55);
			MULT_56(2)<=signed(DIN_56_7)*signed(FMAP_3_56);
			MULT_57(2)<=signed(DIN_57_7)*signed(FMAP_3_57);
			MULT_58(2)<=signed(DIN_58_7)*signed(FMAP_3_58);
			MULT_59(2)<=signed(DIN_59_7)*signed(FMAP_3_59);
			MULT_60(2)<=signed(DIN_60_7)*signed(FMAP_3_60);
			MULT_61(2)<=signed(DIN_61_7)*signed(FMAP_3_61);
			MULT_62(2)<=signed(DIN_62_7)*signed(FMAP_3_62);
			MULT_63(2)<=signed(DIN_63_7)*signed(FMAP_3_63);
			MULT_64(2)<=signed(DIN_64_7)*signed(FMAP_3_64);
			MULT_65(2)<=signed(DIN_65_7)*signed(FMAP_3_65);
			MULT_66(2)<=signed(DIN_66_7)*signed(FMAP_3_66);
			MULT_67(2)<=signed(DIN_67_7)*signed(FMAP_3_67);
			MULT_68(2)<=signed(DIN_68_7)*signed(FMAP_3_68);
			MULT_69(2)<=signed(DIN_69_7)*signed(FMAP_3_69);
			MULT_70(2)<=signed(DIN_70_7)*signed(FMAP_3_70);
			MULT_71(2)<=signed(DIN_71_7)*signed(FMAP_3_71);
			MULT_72(2)<=signed(DIN_72_7)*signed(FMAP_3_72);
			MULT_73(2)<=signed(DIN_73_7)*signed(FMAP_3_73);
			MULT_74(2)<=signed(DIN_74_7)*signed(FMAP_3_74);
			MULT_75(2)<=signed(DIN_75_7)*signed(FMAP_3_75);
			MULT_76(2)<=signed(DIN_76_7)*signed(FMAP_3_76);
			MULT_77(2)<=signed(DIN_77_7)*signed(FMAP_3_77);
			MULT_78(2)<=signed(DIN_78_7)*signed(FMAP_3_78);
			MULT_79(2)<=signed(DIN_79_7)*signed(FMAP_3_79);
			MULT_80(2)<=signed(DIN_80_7)*signed(FMAP_3_80);
			MULT_81(2)<=signed(DIN_81_7)*signed(FMAP_3_81);
			MULT_82(2)<=signed(DIN_82_7)*signed(FMAP_3_82);
			MULT_83(2)<=signed(DIN_83_7)*signed(FMAP_3_83);
			MULT_84(2)<=signed(DIN_84_7)*signed(FMAP_3_84);
			MULT_85(2)<=signed(DIN_85_7)*signed(FMAP_3_85);
			MULT_86(2)<=signed(DIN_86_7)*signed(FMAP_3_86);
			MULT_87(2)<=signed(DIN_87_7)*signed(FMAP_3_87);
			MULT_88(2)<=signed(DIN_88_7)*signed(FMAP_3_88);
			MULT_89(2)<=signed(DIN_89_7)*signed(FMAP_3_89);
			MULT_90(2)<=signed(DIN_90_7)*signed(FMAP_3_90);
			MULT_91(2)<=signed(DIN_91_7)*signed(FMAP_3_91);
			MULT_92(2)<=signed(DIN_92_7)*signed(FMAP_3_92);
			MULT_93(2)<=signed(DIN_93_7)*signed(FMAP_3_93);
			MULT_94(2)<=signed(DIN_94_7)*signed(FMAP_3_94);
			MULT_95(2)<=signed(DIN_95_7)*signed(FMAP_3_95);
			MULT_96(2)<=signed(DIN_96_7)*signed(FMAP_3_96);
			MULT_97(2)<=signed(DIN_97_7)*signed(FMAP_3_97);
			MULT_98(2)<=signed(DIN_98_7)*signed(FMAP_3_98);
			MULT_99(2)<=signed(DIN_99_7)*signed(FMAP_3_99);
			MULT_100(2)<=signed(DIN_100_7)*signed(FMAP_3_100);
			MULT_101(2)<=signed(DIN_101_7)*signed(FMAP_3_101);
			MULT_102(2)<=signed(DIN_102_7)*signed(FMAP_3_102);
			MULT_103(2)<=signed(DIN_103_7)*signed(FMAP_3_103);
			MULT_104(2)<=signed(DIN_104_7)*signed(FMAP_3_104);
			MULT_105(2)<=signed(DIN_105_7)*signed(FMAP_3_105);
			MULT_106(2)<=signed(DIN_106_7)*signed(FMAP_3_106);
			MULT_107(2)<=signed(DIN_107_7)*signed(FMAP_3_107);
			MULT_108(2)<=signed(DIN_108_7)*signed(FMAP_3_108);
			MULT_109(2)<=signed(DIN_109_7)*signed(FMAP_3_109);
			MULT_110(2)<=signed(DIN_110_7)*signed(FMAP_3_110);
			MULT_111(2)<=signed(DIN_111_7)*signed(FMAP_3_111);
			MULT_112(2)<=signed(DIN_112_7)*signed(FMAP_3_112);
			MULT_113(2)<=signed(DIN_113_7)*signed(FMAP_3_113);
			MULT_114(2)<=signed(DIN_114_7)*signed(FMAP_3_114);
			MULT_115(2)<=signed(DIN_115_7)*signed(FMAP_3_115);
			MULT_116(2)<=signed(DIN_116_7)*signed(FMAP_3_116);
			MULT_117(2)<=signed(DIN_117_7)*signed(FMAP_3_117);
			MULT_118(2)<=signed(DIN_118_7)*signed(FMAP_3_118);
			MULT_119(2)<=signed(DIN_119_7)*signed(FMAP_3_119);
			MULT_120(2)<=signed(DIN_120_7)*signed(FMAP_3_120);

			MULT_1(3)<=signed(DIN_1_7)*signed(FMAP_4_1);
			MULT_2(3)<=signed(DIN_2_7)*signed(FMAP_4_2);
			MULT_3(3)<=signed(DIN_3_7)*signed(FMAP_4_3);
			MULT_4(3)<=signed(DIN_4_7)*signed(FMAP_4_4);
			MULT_5(3)<=signed(DIN_5_7)*signed(FMAP_4_5);
			MULT_6(3)<=signed(DIN_6_7)*signed(FMAP_4_6);
			MULT_7(3)<=signed(DIN_7_7)*signed(FMAP_4_7);
			MULT_8(3)<=signed(DIN_8_7)*signed(FMAP_4_8);
			MULT_9(3)<=signed(DIN_9_7)*signed(FMAP_4_9);
			MULT_10(3)<=signed(DIN_10_7)*signed(FMAP_4_10);
			MULT_11(3)<=signed(DIN_11_7)*signed(FMAP_4_11);
			MULT_12(3)<=signed(DIN_12_7)*signed(FMAP_4_12);
			MULT_13(3)<=signed(DIN_13_7)*signed(FMAP_4_13);
			MULT_14(3)<=signed(DIN_14_7)*signed(FMAP_4_14);
			MULT_15(3)<=signed(DIN_15_7)*signed(FMAP_4_15);
			MULT_16(3)<=signed(DIN_16_7)*signed(FMAP_4_16);
			MULT_17(3)<=signed(DIN_17_7)*signed(FMAP_4_17);
			MULT_18(3)<=signed(DIN_18_7)*signed(FMAP_4_18);
			MULT_19(3)<=signed(DIN_19_7)*signed(FMAP_4_19);
			MULT_20(3)<=signed(DIN_20_7)*signed(FMAP_4_20);
			MULT_21(3)<=signed(DIN_21_7)*signed(FMAP_4_21);
			MULT_22(3)<=signed(DIN_22_7)*signed(FMAP_4_22);
			MULT_23(3)<=signed(DIN_23_7)*signed(FMAP_4_23);
			MULT_24(3)<=signed(DIN_24_7)*signed(FMAP_4_24);
			MULT_25(3)<=signed(DIN_25_7)*signed(FMAP_4_25);
			MULT_26(3)<=signed(DIN_26_7)*signed(FMAP_4_26);
			MULT_27(3)<=signed(DIN_27_7)*signed(FMAP_4_27);
			MULT_28(3)<=signed(DIN_28_7)*signed(FMAP_4_28);
			MULT_29(3)<=signed(DIN_29_7)*signed(FMAP_4_29);
			MULT_30(3)<=signed(DIN_30_7)*signed(FMAP_4_30);
			MULT_31(3)<=signed(DIN_31_7)*signed(FMAP_4_31);
			MULT_32(3)<=signed(DIN_32_7)*signed(FMAP_4_32);
			MULT_33(3)<=signed(DIN_33_7)*signed(FMAP_4_33);
			MULT_34(3)<=signed(DIN_34_7)*signed(FMAP_4_34);
			MULT_35(3)<=signed(DIN_35_7)*signed(FMAP_4_35);
			MULT_36(3)<=signed(DIN_36_7)*signed(FMAP_4_36);
			MULT_37(3)<=signed(DIN_37_7)*signed(FMAP_4_37);
			MULT_38(3)<=signed(DIN_38_7)*signed(FMAP_4_38);
			MULT_39(3)<=signed(DIN_39_7)*signed(FMAP_4_39);
			MULT_40(3)<=signed(DIN_40_7)*signed(FMAP_4_40);
			MULT_41(3)<=signed(DIN_41_7)*signed(FMAP_4_41);
			MULT_42(3)<=signed(DIN_42_7)*signed(FMAP_4_42);
			MULT_43(3)<=signed(DIN_43_7)*signed(FMAP_4_43);
			MULT_44(3)<=signed(DIN_44_7)*signed(FMAP_4_44);
			MULT_45(3)<=signed(DIN_45_7)*signed(FMAP_4_45);
			MULT_46(3)<=signed(DIN_46_7)*signed(FMAP_4_46);
			MULT_47(3)<=signed(DIN_47_7)*signed(FMAP_4_47);
			MULT_48(3)<=signed(DIN_48_7)*signed(FMAP_4_48);
			MULT_49(3)<=signed(DIN_49_7)*signed(FMAP_4_49);
			MULT_50(3)<=signed(DIN_50_7)*signed(FMAP_4_50);
			MULT_51(3)<=signed(DIN_51_7)*signed(FMAP_4_51);
			MULT_52(3)<=signed(DIN_52_7)*signed(FMAP_4_52);
			MULT_53(3)<=signed(DIN_53_7)*signed(FMAP_4_53);
			MULT_54(3)<=signed(DIN_54_7)*signed(FMAP_4_54);
			MULT_55(3)<=signed(DIN_55_7)*signed(FMAP_4_55);
			MULT_56(3)<=signed(DIN_56_7)*signed(FMAP_4_56);
			MULT_57(3)<=signed(DIN_57_7)*signed(FMAP_4_57);
			MULT_58(3)<=signed(DIN_58_7)*signed(FMAP_4_58);
			MULT_59(3)<=signed(DIN_59_7)*signed(FMAP_4_59);
			MULT_60(3)<=signed(DIN_60_7)*signed(FMAP_4_60);
			MULT_61(3)<=signed(DIN_61_7)*signed(FMAP_4_61);
			MULT_62(3)<=signed(DIN_62_7)*signed(FMAP_4_62);
			MULT_63(3)<=signed(DIN_63_7)*signed(FMAP_4_63);
			MULT_64(3)<=signed(DIN_64_7)*signed(FMAP_4_64);
			MULT_65(3)<=signed(DIN_65_7)*signed(FMAP_4_65);
			MULT_66(3)<=signed(DIN_66_7)*signed(FMAP_4_66);
			MULT_67(3)<=signed(DIN_67_7)*signed(FMAP_4_67);
			MULT_68(3)<=signed(DIN_68_7)*signed(FMAP_4_68);
			MULT_69(3)<=signed(DIN_69_7)*signed(FMAP_4_69);
			MULT_70(3)<=signed(DIN_70_7)*signed(FMAP_4_70);
			MULT_71(3)<=signed(DIN_71_7)*signed(FMAP_4_71);
			MULT_72(3)<=signed(DIN_72_7)*signed(FMAP_4_72);
			MULT_73(3)<=signed(DIN_73_7)*signed(FMAP_4_73);
			MULT_74(3)<=signed(DIN_74_7)*signed(FMAP_4_74);
			MULT_75(3)<=signed(DIN_75_7)*signed(FMAP_4_75);
			MULT_76(3)<=signed(DIN_76_7)*signed(FMAP_4_76);
			MULT_77(3)<=signed(DIN_77_7)*signed(FMAP_4_77);
			MULT_78(3)<=signed(DIN_78_7)*signed(FMAP_4_78);
			MULT_79(3)<=signed(DIN_79_7)*signed(FMAP_4_79);
			MULT_80(3)<=signed(DIN_80_7)*signed(FMAP_4_80);
			MULT_81(3)<=signed(DIN_81_7)*signed(FMAP_4_81);
			MULT_82(3)<=signed(DIN_82_7)*signed(FMAP_4_82);
			MULT_83(3)<=signed(DIN_83_7)*signed(FMAP_4_83);
			MULT_84(3)<=signed(DIN_84_7)*signed(FMAP_4_84);
			MULT_85(3)<=signed(DIN_85_7)*signed(FMAP_4_85);
			MULT_86(3)<=signed(DIN_86_7)*signed(FMAP_4_86);
			MULT_87(3)<=signed(DIN_87_7)*signed(FMAP_4_87);
			MULT_88(3)<=signed(DIN_88_7)*signed(FMAP_4_88);
			MULT_89(3)<=signed(DIN_89_7)*signed(FMAP_4_89);
			MULT_90(3)<=signed(DIN_90_7)*signed(FMAP_4_90);
			MULT_91(3)<=signed(DIN_91_7)*signed(FMAP_4_91);
			MULT_92(3)<=signed(DIN_92_7)*signed(FMAP_4_92);
			MULT_93(3)<=signed(DIN_93_7)*signed(FMAP_4_93);
			MULT_94(3)<=signed(DIN_94_7)*signed(FMAP_4_94);
			MULT_95(3)<=signed(DIN_95_7)*signed(FMAP_4_95);
			MULT_96(3)<=signed(DIN_96_7)*signed(FMAP_4_96);
			MULT_97(3)<=signed(DIN_97_7)*signed(FMAP_4_97);
			MULT_98(3)<=signed(DIN_98_7)*signed(FMAP_4_98);
			MULT_99(3)<=signed(DIN_99_7)*signed(FMAP_4_99);
			MULT_100(3)<=signed(DIN_100_7)*signed(FMAP_4_100);
			MULT_101(3)<=signed(DIN_101_7)*signed(FMAP_4_101);
			MULT_102(3)<=signed(DIN_102_7)*signed(FMAP_4_102);
			MULT_103(3)<=signed(DIN_103_7)*signed(FMAP_4_103);
			MULT_104(3)<=signed(DIN_104_7)*signed(FMAP_4_104);
			MULT_105(3)<=signed(DIN_105_7)*signed(FMAP_4_105);
			MULT_106(3)<=signed(DIN_106_7)*signed(FMAP_4_106);
			MULT_107(3)<=signed(DIN_107_7)*signed(FMAP_4_107);
			MULT_108(3)<=signed(DIN_108_7)*signed(FMAP_4_108);
			MULT_109(3)<=signed(DIN_109_7)*signed(FMAP_4_109);
			MULT_110(3)<=signed(DIN_110_7)*signed(FMAP_4_110);
			MULT_111(3)<=signed(DIN_111_7)*signed(FMAP_4_111);
			MULT_112(3)<=signed(DIN_112_7)*signed(FMAP_4_112);
			MULT_113(3)<=signed(DIN_113_7)*signed(FMAP_4_113);
			MULT_114(3)<=signed(DIN_114_7)*signed(FMAP_4_114);
			MULT_115(3)<=signed(DIN_115_7)*signed(FMAP_4_115);
			MULT_116(3)<=signed(DIN_116_7)*signed(FMAP_4_116);
			MULT_117(3)<=signed(DIN_117_7)*signed(FMAP_4_117);
			MULT_118(3)<=signed(DIN_118_7)*signed(FMAP_4_118);
			MULT_119(3)<=signed(DIN_119_7)*signed(FMAP_4_119);
			MULT_120(3)<=signed(DIN_120_7)*signed(FMAP_4_120);

			MULT_1(4)<=signed(DIN_1_7)*signed(FMAP_5_1);
			MULT_2(4)<=signed(DIN_2_7)*signed(FMAP_5_2);
			MULT_3(4)<=signed(DIN_3_7)*signed(FMAP_5_3);
			MULT_4(4)<=signed(DIN_4_7)*signed(FMAP_5_4);
			MULT_5(4)<=signed(DIN_5_7)*signed(FMAP_5_5);
			MULT_6(4)<=signed(DIN_6_7)*signed(FMAP_5_6);
			MULT_7(4)<=signed(DIN_7_7)*signed(FMAP_5_7);
			MULT_8(4)<=signed(DIN_8_7)*signed(FMAP_5_8);
			MULT_9(4)<=signed(DIN_9_7)*signed(FMAP_5_9);
			MULT_10(4)<=signed(DIN_10_7)*signed(FMAP_5_10);
			MULT_11(4)<=signed(DIN_11_7)*signed(FMAP_5_11);
			MULT_12(4)<=signed(DIN_12_7)*signed(FMAP_5_12);
			MULT_13(4)<=signed(DIN_13_7)*signed(FMAP_5_13);
			MULT_14(4)<=signed(DIN_14_7)*signed(FMAP_5_14);
			MULT_15(4)<=signed(DIN_15_7)*signed(FMAP_5_15);
			MULT_16(4)<=signed(DIN_16_7)*signed(FMAP_5_16);
			MULT_17(4)<=signed(DIN_17_7)*signed(FMAP_5_17);
			MULT_18(4)<=signed(DIN_18_7)*signed(FMAP_5_18);
			MULT_19(4)<=signed(DIN_19_7)*signed(FMAP_5_19);
			MULT_20(4)<=signed(DIN_20_7)*signed(FMAP_5_20);
			MULT_21(4)<=signed(DIN_21_7)*signed(FMAP_5_21);
			MULT_22(4)<=signed(DIN_22_7)*signed(FMAP_5_22);
			MULT_23(4)<=signed(DIN_23_7)*signed(FMAP_5_23);
			MULT_24(4)<=signed(DIN_24_7)*signed(FMAP_5_24);
			MULT_25(4)<=signed(DIN_25_7)*signed(FMAP_5_25);
			MULT_26(4)<=signed(DIN_26_7)*signed(FMAP_5_26);
			MULT_27(4)<=signed(DIN_27_7)*signed(FMAP_5_27);
			MULT_28(4)<=signed(DIN_28_7)*signed(FMAP_5_28);
			MULT_29(4)<=signed(DIN_29_7)*signed(FMAP_5_29);
			MULT_30(4)<=signed(DIN_30_7)*signed(FMAP_5_30);
			MULT_31(4)<=signed(DIN_31_7)*signed(FMAP_5_31);
			MULT_32(4)<=signed(DIN_32_7)*signed(FMAP_5_32);
			MULT_33(4)<=signed(DIN_33_7)*signed(FMAP_5_33);
			MULT_34(4)<=signed(DIN_34_7)*signed(FMAP_5_34);
			MULT_35(4)<=signed(DIN_35_7)*signed(FMAP_5_35);
			MULT_36(4)<=signed(DIN_36_7)*signed(FMAP_5_36);
			MULT_37(4)<=signed(DIN_37_7)*signed(FMAP_5_37);
			MULT_38(4)<=signed(DIN_38_7)*signed(FMAP_5_38);
			MULT_39(4)<=signed(DIN_39_7)*signed(FMAP_5_39);
			MULT_40(4)<=signed(DIN_40_7)*signed(FMAP_5_40);
			MULT_41(4)<=signed(DIN_41_7)*signed(FMAP_5_41);
			MULT_42(4)<=signed(DIN_42_7)*signed(FMAP_5_42);
			MULT_43(4)<=signed(DIN_43_7)*signed(FMAP_5_43);
			MULT_44(4)<=signed(DIN_44_7)*signed(FMAP_5_44);
			MULT_45(4)<=signed(DIN_45_7)*signed(FMAP_5_45);
			MULT_46(4)<=signed(DIN_46_7)*signed(FMAP_5_46);
			MULT_47(4)<=signed(DIN_47_7)*signed(FMAP_5_47);
			MULT_48(4)<=signed(DIN_48_7)*signed(FMAP_5_48);
			MULT_49(4)<=signed(DIN_49_7)*signed(FMAP_5_49);
			MULT_50(4)<=signed(DIN_50_7)*signed(FMAP_5_50);
			MULT_51(4)<=signed(DIN_51_7)*signed(FMAP_5_51);
			MULT_52(4)<=signed(DIN_52_7)*signed(FMAP_5_52);
			MULT_53(4)<=signed(DIN_53_7)*signed(FMAP_5_53);
			MULT_54(4)<=signed(DIN_54_7)*signed(FMAP_5_54);
			MULT_55(4)<=signed(DIN_55_7)*signed(FMAP_5_55);
			MULT_56(4)<=signed(DIN_56_7)*signed(FMAP_5_56);
			MULT_57(4)<=signed(DIN_57_7)*signed(FMAP_5_57);
			MULT_58(4)<=signed(DIN_58_7)*signed(FMAP_5_58);
			MULT_59(4)<=signed(DIN_59_7)*signed(FMAP_5_59);
			MULT_60(4)<=signed(DIN_60_7)*signed(FMAP_5_60);
			MULT_61(4)<=signed(DIN_61_7)*signed(FMAP_5_61);
			MULT_62(4)<=signed(DIN_62_7)*signed(FMAP_5_62);
			MULT_63(4)<=signed(DIN_63_7)*signed(FMAP_5_63);
			MULT_64(4)<=signed(DIN_64_7)*signed(FMAP_5_64);
			MULT_65(4)<=signed(DIN_65_7)*signed(FMAP_5_65);
			MULT_66(4)<=signed(DIN_66_7)*signed(FMAP_5_66);
			MULT_67(4)<=signed(DIN_67_7)*signed(FMAP_5_67);
			MULT_68(4)<=signed(DIN_68_7)*signed(FMAP_5_68);
			MULT_69(4)<=signed(DIN_69_7)*signed(FMAP_5_69);
			MULT_70(4)<=signed(DIN_70_7)*signed(FMAP_5_70);
			MULT_71(4)<=signed(DIN_71_7)*signed(FMAP_5_71);
			MULT_72(4)<=signed(DIN_72_7)*signed(FMAP_5_72);
			MULT_73(4)<=signed(DIN_73_7)*signed(FMAP_5_73);
			MULT_74(4)<=signed(DIN_74_7)*signed(FMAP_5_74);
			MULT_75(4)<=signed(DIN_75_7)*signed(FMAP_5_75);
			MULT_76(4)<=signed(DIN_76_7)*signed(FMAP_5_76);
			MULT_77(4)<=signed(DIN_77_7)*signed(FMAP_5_77);
			MULT_78(4)<=signed(DIN_78_7)*signed(FMAP_5_78);
			MULT_79(4)<=signed(DIN_79_7)*signed(FMAP_5_79);
			MULT_80(4)<=signed(DIN_80_7)*signed(FMAP_5_80);
			MULT_81(4)<=signed(DIN_81_7)*signed(FMAP_5_81);
			MULT_82(4)<=signed(DIN_82_7)*signed(FMAP_5_82);
			MULT_83(4)<=signed(DIN_83_7)*signed(FMAP_5_83);
			MULT_84(4)<=signed(DIN_84_7)*signed(FMAP_5_84);
			MULT_85(4)<=signed(DIN_85_7)*signed(FMAP_5_85);
			MULT_86(4)<=signed(DIN_86_7)*signed(FMAP_5_86);
			MULT_87(4)<=signed(DIN_87_7)*signed(FMAP_5_87);
			MULT_88(4)<=signed(DIN_88_7)*signed(FMAP_5_88);
			MULT_89(4)<=signed(DIN_89_7)*signed(FMAP_5_89);
			MULT_90(4)<=signed(DIN_90_7)*signed(FMAP_5_90);
			MULT_91(4)<=signed(DIN_91_7)*signed(FMAP_5_91);
			MULT_92(4)<=signed(DIN_92_7)*signed(FMAP_5_92);
			MULT_93(4)<=signed(DIN_93_7)*signed(FMAP_5_93);
			MULT_94(4)<=signed(DIN_94_7)*signed(FMAP_5_94);
			MULT_95(4)<=signed(DIN_95_7)*signed(FMAP_5_95);
			MULT_96(4)<=signed(DIN_96_7)*signed(FMAP_5_96);
			MULT_97(4)<=signed(DIN_97_7)*signed(FMAP_5_97);
			MULT_98(4)<=signed(DIN_98_7)*signed(FMAP_5_98);
			MULT_99(4)<=signed(DIN_99_7)*signed(FMAP_5_99);
			MULT_100(4)<=signed(DIN_100_7)*signed(FMAP_5_100);
			MULT_101(4)<=signed(DIN_101_7)*signed(FMAP_5_101);
			MULT_102(4)<=signed(DIN_102_7)*signed(FMAP_5_102);
			MULT_103(4)<=signed(DIN_103_7)*signed(FMAP_5_103);
			MULT_104(4)<=signed(DIN_104_7)*signed(FMAP_5_104);
			MULT_105(4)<=signed(DIN_105_7)*signed(FMAP_5_105);
			MULT_106(4)<=signed(DIN_106_7)*signed(FMAP_5_106);
			MULT_107(4)<=signed(DIN_107_7)*signed(FMAP_5_107);
			MULT_108(4)<=signed(DIN_108_7)*signed(FMAP_5_108);
			MULT_109(4)<=signed(DIN_109_7)*signed(FMAP_5_109);
			MULT_110(4)<=signed(DIN_110_7)*signed(FMAP_5_110);
			MULT_111(4)<=signed(DIN_111_7)*signed(FMAP_5_111);
			MULT_112(4)<=signed(DIN_112_7)*signed(FMAP_5_112);
			MULT_113(4)<=signed(DIN_113_7)*signed(FMAP_5_113);
			MULT_114(4)<=signed(DIN_114_7)*signed(FMAP_5_114);
			MULT_115(4)<=signed(DIN_115_7)*signed(FMAP_5_115);
			MULT_116(4)<=signed(DIN_116_7)*signed(FMAP_5_116);
			MULT_117(4)<=signed(DIN_117_7)*signed(FMAP_5_117);
			MULT_118(4)<=signed(DIN_118_7)*signed(FMAP_5_118);
			MULT_119(4)<=signed(DIN_119_7)*signed(FMAP_5_119);
			MULT_120(4)<=signed(DIN_120_7)*signed(FMAP_5_120);

			MULT_1(5)<=signed(DIN_1_7)*signed(FMAP_6_1);
			MULT_2(5)<=signed(DIN_2_7)*signed(FMAP_6_2);
			MULT_3(5)<=signed(DIN_3_7)*signed(FMAP_6_3);
			MULT_4(5)<=signed(DIN_4_7)*signed(FMAP_6_4);
			MULT_5(5)<=signed(DIN_5_7)*signed(FMAP_6_5);
			MULT_6(5)<=signed(DIN_6_7)*signed(FMAP_6_6);
			MULT_7(5)<=signed(DIN_7_7)*signed(FMAP_6_7);
			MULT_8(5)<=signed(DIN_8_7)*signed(FMAP_6_8);
			MULT_9(5)<=signed(DIN_9_7)*signed(FMAP_6_9);
			MULT_10(5)<=signed(DIN_10_7)*signed(FMAP_6_10);
			MULT_11(5)<=signed(DIN_11_7)*signed(FMAP_6_11);
			MULT_12(5)<=signed(DIN_12_7)*signed(FMAP_6_12);
			MULT_13(5)<=signed(DIN_13_7)*signed(FMAP_6_13);
			MULT_14(5)<=signed(DIN_14_7)*signed(FMAP_6_14);
			MULT_15(5)<=signed(DIN_15_7)*signed(FMAP_6_15);
			MULT_16(5)<=signed(DIN_16_7)*signed(FMAP_6_16);
			MULT_17(5)<=signed(DIN_17_7)*signed(FMAP_6_17);
			MULT_18(5)<=signed(DIN_18_7)*signed(FMAP_6_18);
			MULT_19(5)<=signed(DIN_19_7)*signed(FMAP_6_19);
			MULT_20(5)<=signed(DIN_20_7)*signed(FMAP_6_20);
			MULT_21(5)<=signed(DIN_21_7)*signed(FMAP_6_21);
			MULT_22(5)<=signed(DIN_22_7)*signed(FMAP_6_22);
			MULT_23(5)<=signed(DIN_23_7)*signed(FMAP_6_23);
			MULT_24(5)<=signed(DIN_24_7)*signed(FMAP_6_24);
			MULT_25(5)<=signed(DIN_25_7)*signed(FMAP_6_25);
			MULT_26(5)<=signed(DIN_26_7)*signed(FMAP_6_26);
			MULT_27(5)<=signed(DIN_27_7)*signed(FMAP_6_27);
			MULT_28(5)<=signed(DIN_28_7)*signed(FMAP_6_28);
			MULT_29(5)<=signed(DIN_29_7)*signed(FMAP_6_29);
			MULT_30(5)<=signed(DIN_30_7)*signed(FMAP_6_30);
			MULT_31(5)<=signed(DIN_31_7)*signed(FMAP_6_31);
			MULT_32(5)<=signed(DIN_32_7)*signed(FMAP_6_32);
			MULT_33(5)<=signed(DIN_33_7)*signed(FMAP_6_33);
			MULT_34(5)<=signed(DIN_34_7)*signed(FMAP_6_34);
			MULT_35(5)<=signed(DIN_35_7)*signed(FMAP_6_35);
			MULT_36(5)<=signed(DIN_36_7)*signed(FMAP_6_36);
			MULT_37(5)<=signed(DIN_37_7)*signed(FMAP_6_37);
			MULT_38(5)<=signed(DIN_38_7)*signed(FMAP_6_38);
			MULT_39(5)<=signed(DIN_39_7)*signed(FMAP_6_39);
			MULT_40(5)<=signed(DIN_40_7)*signed(FMAP_6_40);
			MULT_41(5)<=signed(DIN_41_7)*signed(FMAP_6_41);
			MULT_42(5)<=signed(DIN_42_7)*signed(FMAP_6_42);
			MULT_43(5)<=signed(DIN_43_7)*signed(FMAP_6_43);
			MULT_44(5)<=signed(DIN_44_7)*signed(FMAP_6_44);
			MULT_45(5)<=signed(DIN_45_7)*signed(FMAP_6_45);
			MULT_46(5)<=signed(DIN_46_7)*signed(FMAP_6_46);
			MULT_47(5)<=signed(DIN_47_7)*signed(FMAP_6_47);
			MULT_48(5)<=signed(DIN_48_7)*signed(FMAP_6_48);
			MULT_49(5)<=signed(DIN_49_7)*signed(FMAP_6_49);
			MULT_50(5)<=signed(DIN_50_7)*signed(FMAP_6_50);
			MULT_51(5)<=signed(DIN_51_7)*signed(FMAP_6_51);
			MULT_52(5)<=signed(DIN_52_7)*signed(FMAP_6_52);
			MULT_53(5)<=signed(DIN_53_7)*signed(FMAP_6_53);
			MULT_54(5)<=signed(DIN_54_7)*signed(FMAP_6_54);
			MULT_55(5)<=signed(DIN_55_7)*signed(FMAP_6_55);
			MULT_56(5)<=signed(DIN_56_7)*signed(FMAP_6_56);
			MULT_57(5)<=signed(DIN_57_7)*signed(FMAP_6_57);
			MULT_58(5)<=signed(DIN_58_7)*signed(FMAP_6_58);
			MULT_59(5)<=signed(DIN_59_7)*signed(FMAP_6_59);
			MULT_60(5)<=signed(DIN_60_7)*signed(FMAP_6_60);
			MULT_61(5)<=signed(DIN_61_7)*signed(FMAP_6_61);
			MULT_62(5)<=signed(DIN_62_7)*signed(FMAP_6_62);
			MULT_63(5)<=signed(DIN_63_7)*signed(FMAP_6_63);
			MULT_64(5)<=signed(DIN_64_7)*signed(FMAP_6_64);
			MULT_65(5)<=signed(DIN_65_7)*signed(FMAP_6_65);
			MULT_66(5)<=signed(DIN_66_7)*signed(FMAP_6_66);
			MULT_67(5)<=signed(DIN_67_7)*signed(FMAP_6_67);
			MULT_68(5)<=signed(DIN_68_7)*signed(FMAP_6_68);
			MULT_69(5)<=signed(DIN_69_7)*signed(FMAP_6_69);
			MULT_70(5)<=signed(DIN_70_7)*signed(FMAP_6_70);
			MULT_71(5)<=signed(DIN_71_7)*signed(FMAP_6_71);
			MULT_72(5)<=signed(DIN_72_7)*signed(FMAP_6_72);
			MULT_73(5)<=signed(DIN_73_7)*signed(FMAP_6_73);
			MULT_74(5)<=signed(DIN_74_7)*signed(FMAP_6_74);
			MULT_75(5)<=signed(DIN_75_7)*signed(FMAP_6_75);
			MULT_76(5)<=signed(DIN_76_7)*signed(FMAP_6_76);
			MULT_77(5)<=signed(DIN_77_7)*signed(FMAP_6_77);
			MULT_78(5)<=signed(DIN_78_7)*signed(FMAP_6_78);
			MULT_79(5)<=signed(DIN_79_7)*signed(FMAP_6_79);
			MULT_80(5)<=signed(DIN_80_7)*signed(FMAP_6_80);
			MULT_81(5)<=signed(DIN_81_7)*signed(FMAP_6_81);
			MULT_82(5)<=signed(DIN_82_7)*signed(FMAP_6_82);
			MULT_83(5)<=signed(DIN_83_7)*signed(FMAP_6_83);
			MULT_84(5)<=signed(DIN_84_7)*signed(FMAP_6_84);
			MULT_85(5)<=signed(DIN_85_7)*signed(FMAP_6_85);
			MULT_86(5)<=signed(DIN_86_7)*signed(FMAP_6_86);
			MULT_87(5)<=signed(DIN_87_7)*signed(FMAP_6_87);
			MULT_88(5)<=signed(DIN_88_7)*signed(FMAP_6_88);
			MULT_89(5)<=signed(DIN_89_7)*signed(FMAP_6_89);
			MULT_90(5)<=signed(DIN_90_7)*signed(FMAP_6_90);
			MULT_91(5)<=signed(DIN_91_7)*signed(FMAP_6_91);
			MULT_92(5)<=signed(DIN_92_7)*signed(FMAP_6_92);
			MULT_93(5)<=signed(DIN_93_7)*signed(FMAP_6_93);
			MULT_94(5)<=signed(DIN_94_7)*signed(FMAP_6_94);
			MULT_95(5)<=signed(DIN_95_7)*signed(FMAP_6_95);
			MULT_96(5)<=signed(DIN_96_7)*signed(FMAP_6_96);
			MULT_97(5)<=signed(DIN_97_7)*signed(FMAP_6_97);
			MULT_98(5)<=signed(DIN_98_7)*signed(FMAP_6_98);
			MULT_99(5)<=signed(DIN_99_7)*signed(FMAP_6_99);
			MULT_100(5)<=signed(DIN_100_7)*signed(FMAP_6_100);
			MULT_101(5)<=signed(DIN_101_7)*signed(FMAP_6_101);
			MULT_102(5)<=signed(DIN_102_7)*signed(FMAP_6_102);
			MULT_103(5)<=signed(DIN_103_7)*signed(FMAP_6_103);
			MULT_104(5)<=signed(DIN_104_7)*signed(FMAP_6_104);
			MULT_105(5)<=signed(DIN_105_7)*signed(FMAP_6_105);
			MULT_106(5)<=signed(DIN_106_7)*signed(FMAP_6_106);
			MULT_107(5)<=signed(DIN_107_7)*signed(FMAP_6_107);
			MULT_108(5)<=signed(DIN_108_7)*signed(FMAP_6_108);
			MULT_109(5)<=signed(DIN_109_7)*signed(FMAP_6_109);
			MULT_110(5)<=signed(DIN_110_7)*signed(FMAP_6_110);
			MULT_111(5)<=signed(DIN_111_7)*signed(FMAP_6_111);
			MULT_112(5)<=signed(DIN_112_7)*signed(FMAP_6_112);
			MULT_113(5)<=signed(DIN_113_7)*signed(FMAP_6_113);
			MULT_114(5)<=signed(DIN_114_7)*signed(FMAP_6_114);
			MULT_115(5)<=signed(DIN_115_7)*signed(FMAP_6_115);
			MULT_116(5)<=signed(DIN_116_7)*signed(FMAP_6_116);
			MULT_117(5)<=signed(DIN_117_7)*signed(FMAP_6_117);
			MULT_118(5)<=signed(DIN_118_7)*signed(FMAP_6_118);
			MULT_119(5)<=signed(DIN_119_7)*signed(FMAP_6_119);
			MULT_120(5)<=signed(DIN_120_7)*signed(FMAP_6_120);

			MULT_1(6)<=signed(DIN_1_7)*signed(FMAP_7_1);
			MULT_2(6)<=signed(DIN_2_7)*signed(FMAP_7_2);
			MULT_3(6)<=signed(DIN_3_7)*signed(FMAP_7_3);
			MULT_4(6)<=signed(DIN_4_7)*signed(FMAP_7_4);
			MULT_5(6)<=signed(DIN_5_7)*signed(FMAP_7_5);
			MULT_6(6)<=signed(DIN_6_7)*signed(FMAP_7_6);
			MULT_7(6)<=signed(DIN_7_7)*signed(FMAP_7_7);
			MULT_8(6)<=signed(DIN_8_7)*signed(FMAP_7_8);
			MULT_9(6)<=signed(DIN_9_7)*signed(FMAP_7_9);
			MULT_10(6)<=signed(DIN_10_7)*signed(FMAP_7_10);
			MULT_11(6)<=signed(DIN_11_7)*signed(FMAP_7_11);
			MULT_12(6)<=signed(DIN_12_7)*signed(FMAP_7_12);
			MULT_13(6)<=signed(DIN_13_7)*signed(FMAP_7_13);
			MULT_14(6)<=signed(DIN_14_7)*signed(FMAP_7_14);
			MULT_15(6)<=signed(DIN_15_7)*signed(FMAP_7_15);
			MULT_16(6)<=signed(DIN_16_7)*signed(FMAP_7_16);
			MULT_17(6)<=signed(DIN_17_7)*signed(FMAP_7_17);
			MULT_18(6)<=signed(DIN_18_7)*signed(FMAP_7_18);
			MULT_19(6)<=signed(DIN_19_7)*signed(FMAP_7_19);
			MULT_20(6)<=signed(DIN_20_7)*signed(FMAP_7_20);
			MULT_21(6)<=signed(DIN_21_7)*signed(FMAP_7_21);
			MULT_22(6)<=signed(DIN_22_7)*signed(FMAP_7_22);
			MULT_23(6)<=signed(DIN_23_7)*signed(FMAP_7_23);
			MULT_24(6)<=signed(DIN_24_7)*signed(FMAP_7_24);
			MULT_25(6)<=signed(DIN_25_7)*signed(FMAP_7_25);
			MULT_26(6)<=signed(DIN_26_7)*signed(FMAP_7_26);
			MULT_27(6)<=signed(DIN_27_7)*signed(FMAP_7_27);
			MULT_28(6)<=signed(DIN_28_7)*signed(FMAP_7_28);
			MULT_29(6)<=signed(DIN_29_7)*signed(FMAP_7_29);
			MULT_30(6)<=signed(DIN_30_7)*signed(FMAP_7_30);
			MULT_31(6)<=signed(DIN_31_7)*signed(FMAP_7_31);
			MULT_32(6)<=signed(DIN_32_7)*signed(FMAP_7_32);
			MULT_33(6)<=signed(DIN_33_7)*signed(FMAP_7_33);
			MULT_34(6)<=signed(DIN_34_7)*signed(FMAP_7_34);
			MULT_35(6)<=signed(DIN_35_7)*signed(FMAP_7_35);
			MULT_36(6)<=signed(DIN_36_7)*signed(FMAP_7_36);
			MULT_37(6)<=signed(DIN_37_7)*signed(FMAP_7_37);
			MULT_38(6)<=signed(DIN_38_7)*signed(FMAP_7_38);
			MULT_39(6)<=signed(DIN_39_7)*signed(FMAP_7_39);
			MULT_40(6)<=signed(DIN_40_7)*signed(FMAP_7_40);
			MULT_41(6)<=signed(DIN_41_7)*signed(FMAP_7_41);
			MULT_42(6)<=signed(DIN_42_7)*signed(FMAP_7_42);
			MULT_43(6)<=signed(DIN_43_7)*signed(FMAP_7_43);
			MULT_44(6)<=signed(DIN_44_7)*signed(FMAP_7_44);
			MULT_45(6)<=signed(DIN_45_7)*signed(FMAP_7_45);
			MULT_46(6)<=signed(DIN_46_7)*signed(FMAP_7_46);
			MULT_47(6)<=signed(DIN_47_7)*signed(FMAP_7_47);
			MULT_48(6)<=signed(DIN_48_7)*signed(FMAP_7_48);
			MULT_49(6)<=signed(DIN_49_7)*signed(FMAP_7_49);
			MULT_50(6)<=signed(DIN_50_7)*signed(FMAP_7_50);
			MULT_51(6)<=signed(DIN_51_7)*signed(FMAP_7_51);
			MULT_52(6)<=signed(DIN_52_7)*signed(FMAP_7_52);
			MULT_53(6)<=signed(DIN_53_7)*signed(FMAP_7_53);
			MULT_54(6)<=signed(DIN_54_7)*signed(FMAP_7_54);
			MULT_55(6)<=signed(DIN_55_7)*signed(FMAP_7_55);
			MULT_56(6)<=signed(DIN_56_7)*signed(FMAP_7_56);
			MULT_57(6)<=signed(DIN_57_7)*signed(FMAP_7_57);
			MULT_58(6)<=signed(DIN_58_7)*signed(FMAP_7_58);
			MULT_59(6)<=signed(DIN_59_7)*signed(FMAP_7_59);
			MULT_60(6)<=signed(DIN_60_7)*signed(FMAP_7_60);
			MULT_61(6)<=signed(DIN_61_7)*signed(FMAP_7_61);
			MULT_62(6)<=signed(DIN_62_7)*signed(FMAP_7_62);
			MULT_63(6)<=signed(DIN_63_7)*signed(FMAP_7_63);
			MULT_64(6)<=signed(DIN_64_7)*signed(FMAP_7_64);
			MULT_65(6)<=signed(DIN_65_7)*signed(FMAP_7_65);
			MULT_66(6)<=signed(DIN_66_7)*signed(FMAP_7_66);
			MULT_67(6)<=signed(DIN_67_7)*signed(FMAP_7_67);
			MULT_68(6)<=signed(DIN_68_7)*signed(FMAP_7_68);
			MULT_69(6)<=signed(DIN_69_7)*signed(FMAP_7_69);
			MULT_70(6)<=signed(DIN_70_7)*signed(FMAP_7_70);
			MULT_71(6)<=signed(DIN_71_7)*signed(FMAP_7_71);
			MULT_72(6)<=signed(DIN_72_7)*signed(FMAP_7_72);
			MULT_73(6)<=signed(DIN_73_7)*signed(FMAP_7_73);
			MULT_74(6)<=signed(DIN_74_7)*signed(FMAP_7_74);
			MULT_75(6)<=signed(DIN_75_7)*signed(FMAP_7_75);
			MULT_76(6)<=signed(DIN_76_7)*signed(FMAP_7_76);
			MULT_77(6)<=signed(DIN_77_7)*signed(FMAP_7_77);
			MULT_78(6)<=signed(DIN_78_7)*signed(FMAP_7_78);
			MULT_79(6)<=signed(DIN_79_7)*signed(FMAP_7_79);
			MULT_80(6)<=signed(DIN_80_7)*signed(FMAP_7_80);
			MULT_81(6)<=signed(DIN_81_7)*signed(FMAP_7_81);
			MULT_82(6)<=signed(DIN_82_7)*signed(FMAP_7_82);
			MULT_83(6)<=signed(DIN_83_7)*signed(FMAP_7_83);
			MULT_84(6)<=signed(DIN_84_7)*signed(FMAP_7_84);
			MULT_85(6)<=signed(DIN_85_7)*signed(FMAP_7_85);
			MULT_86(6)<=signed(DIN_86_7)*signed(FMAP_7_86);
			MULT_87(6)<=signed(DIN_87_7)*signed(FMAP_7_87);
			MULT_88(6)<=signed(DIN_88_7)*signed(FMAP_7_88);
			MULT_89(6)<=signed(DIN_89_7)*signed(FMAP_7_89);
			MULT_90(6)<=signed(DIN_90_7)*signed(FMAP_7_90);
			MULT_91(6)<=signed(DIN_91_7)*signed(FMAP_7_91);
			MULT_92(6)<=signed(DIN_92_7)*signed(FMAP_7_92);
			MULT_93(6)<=signed(DIN_93_7)*signed(FMAP_7_93);
			MULT_94(6)<=signed(DIN_94_7)*signed(FMAP_7_94);
			MULT_95(6)<=signed(DIN_95_7)*signed(FMAP_7_95);
			MULT_96(6)<=signed(DIN_96_7)*signed(FMAP_7_96);
			MULT_97(6)<=signed(DIN_97_7)*signed(FMAP_7_97);
			MULT_98(6)<=signed(DIN_98_7)*signed(FMAP_7_98);
			MULT_99(6)<=signed(DIN_99_7)*signed(FMAP_7_99);
			MULT_100(6)<=signed(DIN_100_7)*signed(FMAP_7_100);
			MULT_101(6)<=signed(DIN_101_7)*signed(FMAP_7_101);
			MULT_102(6)<=signed(DIN_102_7)*signed(FMAP_7_102);
			MULT_103(6)<=signed(DIN_103_7)*signed(FMAP_7_103);
			MULT_104(6)<=signed(DIN_104_7)*signed(FMAP_7_104);
			MULT_105(6)<=signed(DIN_105_7)*signed(FMAP_7_105);
			MULT_106(6)<=signed(DIN_106_7)*signed(FMAP_7_106);
			MULT_107(6)<=signed(DIN_107_7)*signed(FMAP_7_107);
			MULT_108(6)<=signed(DIN_108_7)*signed(FMAP_7_108);
			MULT_109(6)<=signed(DIN_109_7)*signed(FMAP_7_109);
			MULT_110(6)<=signed(DIN_110_7)*signed(FMAP_7_110);
			MULT_111(6)<=signed(DIN_111_7)*signed(FMAP_7_111);
			MULT_112(6)<=signed(DIN_112_7)*signed(FMAP_7_112);
			MULT_113(6)<=signed(DIN_113_7)*signed(FMAP_7_113);
			MULT_114(6)<=signed(DIN_114_7)*signed(FMAP_7_114);
			MULT_115(6)<=signed(DIN_115_7)*signed(FMAP_7_115);
			MULT_116(6)<=signed(DIN_116_7)*signed(FMAP_7_116);
			MULT_117(6)<=signed(DIN_117_7)*signed(FMAP_7_117);
			MULT_118(6)<=signed(DIN_118_7)*signed(FMAP_7_118);
			MULT_119(6)<=signed(DIN_119_7)*signed(FMAP_7_119);
			MULT_120(6)<=signed(DIN_120_7)*signed(FMAP_7_120);

			MULT_1(7)<=signed(DIN_1_7)*signed(FMAP_8_1);
			MULT_2(7)<=signed(DIN_2_7)*signed(FMAP_8_2);
			MULT_3(7)<=signed(DIN_3_7)*signed(FMAP_8_3);
			MULT_4(7)<=signed(DIN_4_7)*signed(FMAP_8_4);
			MULT_5(7)<=signed(DIN_5_7)*signed(FMAP_8_5);
			MULT_6(7)<=signed(DIN_6_7)*signed(FMAP_8_6);
			MULT_7(7)<=signed(DIN_7_7)*signed(FMAP_8_7);
			MULT_8(7)<=signed(DIN_8_7)*signed(FMAP_8_8);
			MULT_9(7)<=signed(DIN_9_7)*signed(FMAP_8_9);
			MULT_10(7)<=signed(DIN_10_7)*signed(FMAP_8_10);
			MULT_11(7)<=signed(DIN_11_7)*signed(FMAP_8_11);
			MULT_12(7)<=signed(DIN_12_7)*signed(FMAP_8_12);
			MULT_13(7)<=signed(DIN_13_7)*signed(FMAP_8_13);
			MULT_14(7)<=signed(DIN_14_7)*signed(FMAP_8_14);
			MULT_15(7)<=signed(DIN_15_7)*signed(FMAP_8_15);
			MULT_16(7)<=signed(DIN_16_7)*signed(FMAP_8_16);
			MULT_17(7)<=signed(DIN_17_7)*signed(FMAP_8_17);
			MULT_18(7)<=signed(DIN_18_7)*signed(FMAP_8_18);
			MULT_19(7)<=signed(DIN_19_7)*signed(FMAP_8_19);
			MULT_20(7)<=signed(DIN_20_7)*signed(FMAP_8_20);
			MULT_21(7)<=signed(DIN_21_7)*signed(FMAP_8_21);
			MULT_22(7)<=signed(DIN_22_7)*signed(FMAP_8_22);
			MULT_23(7)<=signed(DIN_23_7)*signed(FMAP_8_23);
			MULT_24(7)<=signed(DIN_24_7)*signed(FMAP_8_24);
			MULT_25(7)<=signed(DIN_25_7)*signed(FMAP_8_25);
			MULT_26(7)<=signed(DIN_26_7)*signed(FMAP_8_26);
			MULT_27(7)<=signed(DIN_27_7)*signed(FMAP_8_27);
			MULT_28(7)<=signed(DIN_28_7)*signed(FMAP_8_28);
			MULT_29(7)<=signed(DIN_29_7)*signed(FMAP_8_29);
			MULT_30(7)<=signed(DIN_30_7)*signed(FMAP_8_30);
			MULT_31(7)<=signed(DIN_31_7)*signed(FMAP_8_31);
			MULT_32(7)<=signed(DIN_32_7)*signed(FMAP_8_32);
			MULT_33(7)<=signed(DIN_33_7)*signed(FMAP_8_33);
			MULT_34(7)<=signed(DIN_34_7)*signed(FMAP_8_34);
			MULT_35(7)<=signed(DIN_35_7)*signed(FMAP_8_35);
			MULT_36(7)<=signed(DIN_36_7)*signed(FMAP_8_36);
			MULT_37(7)<=signed(DIN_37_7)*signed(FMAP_8_37);
			MULT_38(7)<=signed(DIN_38_7)*signed(FMAP_8_38);
			MULT_39(7)<=signed(DIN_39_7)*signed(FMAP_8_39);
			MULT_40(7)<=signed(DIN_40_7)*signed(FMAP_8_40);
			MULT_41(7)<=signed(DIN_41_7)*signed(FMAP_8_41);
			MULT_42(7)<=signed(DIN_42_7)*signed(FMAP_8_42);
			MULT_43(7)<=signed(DIN_43_7)*signed(FMAP_8_43);
			MULT_44(7)<=signed(DIN_44_7)*signed(FMAP_8_44);
			MULT_45(7)<=signed(DIN_45_7)*signed(FMAP_8_45);
			MULT_46(7)<=signed(DIN_46_7)*signed(FMAP_8_46);
			MULT_47(7)<=signed(DIN_47_7)*signed(FMAP_8_47);
			MULT_48(7)<=signed(DIN_48_7)*signed(FMAP_8_48);
			MULT_49(7)<=signed(DIN_49_7)*signed(FMAP_8_49);
			MULT_50(7)<=signed(DIN_50_7)*signed(FMAP_8_50);
			MULT_51(7)<=signed(DIN_51_7)*signed(FMAP_8_51);
			MULT_52(7)<=signed(DIN_52_7)*signed(FMAP_8_52);
			MULT_53(7)<=signed(DIN_53_7)*signed(FMAP_8_53);
			MULT_54(7)<=signed(DIN_54_7)*signed(FMAP_8_54);
			MULT_55(7)<=signed(DIN_55_7)*signed(FMAP_8_55);
			MULT_56(7)<=signed(DIN_56_7)*signed(FMAP_8_56);
			MULT_57(7)<=signed(DIN_57_7)*signed(FMAP_8_57);
			MULT_58(7)<=signed(DIN_58_7)*signed(FMAP_8_58);
			MULT_59(7)<=signed(DIN_59_7)*signed(FMAP_8_59);
			MULT_60(7)<=signed(DIN_60_7)*signed(FMAP_8_60);
			MULT_61(7)<=signed(DIN_61_7)*signed(FMAP_8_61);
			MULT_62(7)<=signed(DIN_62_7)*signed(FMAP_8_62);
			MULT_63(7)<=signed(DIN_63_7)*signed(FMAP_8_63);
			MULT_64(7)<=signed(DIN_64_7)*signed(FMAP_8_64);
			MULT_65(7)<=signed(DIN_65_7)*signed(FMAP_8_65);
			MULT_66(7)<=signed(DIN_66_7)*signed(FMAP_8_66);
			MULT_67(7)<=signed(DIN_67_7)*signed(FMAP_8_67);
			MULT_68(7)<=signed(DIN_68_7)*signed(FMAP_8_68);
			MULT_69(7)<=signed(DIN_69_7)*signed(FMAP_8_69);
			MULT_70(7)<=signed(DIN_70_7)*signed(FMAP_8_70);
			MULT_71(7)<=signed(DIN_71_7)*signed(FMAP_8_71);
			MULT_72(7)<=signed(DIN_72_7)*signed(FMAP_8_72);
			MULT_73(7)<=signed(DIN_73_7)*signed(FMAP_8_73);
			MULT_74(7)<=signed(DIN_74_7)*signed(FMAP_8_74);
			MULT_75(7)<=signed(DIN_75_7)*signed(FMAP_8_75);
			MULT_76(7)<=signed(DIN_76_7)*signed(FMAP_8_76);
			MULT_77(7)<=signed(DIN_77_7)*signed(FMAP_8_77);
			MULT_78(7)<=signed(DIN_78_7)*signed(FMAP_8_78);
			MULT_79(7)<=signed(DIN_79_7)*signed(FMAP_8_79);
			MULT_80(7)<=signed(DIN_80_7)*signed(FMAP_8_80);
			MULT_81(7)<=signed(DIN_81_7)*signed(FMAP_8_81);
			MULT_82(7)<=signed(DIN_82_7)*signed(FMAP_8_82);
			MULT_83(7)<=signed(DIN_83_7)*signed(FMAP_8_83);
			MULT_84(7)<=signed(DIN_84_7)*signed(FMAP_8_84);
			MULT_85(7)<=signed(DIN_85_7)*signed(FMAP_8_85);
			MULT_86(7)<=signed(DIN_86_7)*signed(FMAP_8_86);
			MULT_87(7)<=signed(DIN_87_7)*signed(FMAP_8_87);
			MULT_88(7)<=signed(DIN_88_7)*signed(FMAP_8_88);
			MULT_89(7)<=signed(DIN_89_7)*signed(FMAP_8_89);
			MULT_90(7)<=signed(DIN_90_7)*signed(FMAP_8_90);
			MULT_91(7)<=signed(DIN_91_7)*signed(FMAP_8_91);
			MULT_92(7)<=signed(DIN_92_7)*signed(FMAP_8_92);
			MULT_93(7)<=signed(DIN_93_7)*signed(FMAP_8_93);
			MULT_94(7)<=signed(DIN_94_7)*signed(FMAP_8_94);
			MULT_95(7)<=signed(DIN_95_7)*signed(FMAP_8_95);
			MULT_96(7)<=signed(DIN_96_7)*signed(FMAP_8_96);
			MULT_97(7)<=signed(DIN_97_7)*signed(FMAP_8_97);
			MULT_98(7)<=signed(DIN_98_7)*signed(FMAP_8_98);
			MULT_99(7)<=signed(DIN_99_7)*signed(FMAP_8_99);
			MULT_100(7)<=signed(DIN_100_7)*signed(FMAP_8_100);
			MULT_101(7)<=signed(DIN_101_7)*signed(FMAP_8_101);
			MULT_102(7)<=signed(DIN_102_7)*signed(FMAP_8_102);
			MULT_103(7)<=signed(DIN_103_7)*signed(FMAP_8_103);
			MULT_104(7)<=signed(DIN_104_7)*signed(FMAP_8_104);
			MULT_105(7)<=signed(DIN_105_7)*signed(FMAP_8_105);
			MULT_106(7)<=signed(DIN_106_7)*signed(FMAP_8_106);
			MULT_107(7)<=signed(DIN_107_7)*signed(FMAP_8_107);
			MULT_108(7)<=signed(DIN_108_7)*signed(FMAP_8_108);
			MULT_109(7)<=signed(DIN_109_7)*signed(FMAP_8_109);
			MULT_110(7)<=signed(DIN_110_7)*signed(FMAP_8_110);
			MULT_111(7)<=signed(DIN_111_7)*signed(FMAP_8_111);
			MULT_112(7)<=signed(DIN_112_7)*signed(FMAP_8_112);
			MULT_113(7)<=signed(DIN_113_7)*signed(FMAP_8_113);
			MULT_114(7)<=signed(DIN_114_7)*signed(FMAP_8_114);
			MULT_115(7)<=signed(DIN_115_7)*signed(FMAP_8_115);
			MULT_116(7)<=signed(DIN_116_7)*signed(FMAP_8_116);
			MULT_117(7)<=signed(DIN_117_7)*signed(FMAP_8_117);
			MULT_118(7)<=signed(DIN_118_7)*signed(FMAP_8_118);
			MULT_119(7)<=signed(DIN_119_7)*signed(FMAP_8_119);
			MULT_120(7)<=signed(DIN_120_7)*signed(FMAP_8_120);

			MULT_1(8)<=signed(DIN_1_7)*signed(FMAP_9_1);
			MULT_2(8)<=signed(DIN_2_7)*signed(FMAP_9_2);
			MULT_3(8)<=signed(DIN_3_7)*signed(FMAP_9_3);
			MULT_4(8)<=signed(DIN_4_7)*signed(FMAP_9_4);
			MULT_5(8)<=signed(DIN_5_7)*signed(FMAP_9_5);
			MULT_6(8)<=signed(DIN_6_7)*signed(FMAP_9_6);
			MULT_7(8)<=signed(DIN_7_7)*signed(FMAP_9_7);
			MULT_8(8)<=signed(DIN_8_7)*signed(FMAP_9_8);
			MULT_9(8)<=signed(DIN_9_7)*signed(FMAP_9_9);
			MULT_10(8)<=signed(DIN_10_7)*signed(FMAP_9_10);
			MULT_11(8)<=signed(DIN_11_7)*signed(FMAP_9_11);
			MULT_12(8)<=signed(DIN_12_7)*signed(FMAP_9_12);
			MULT_13(8)<=signed(DIN_13_7)*signed(FMAP_9_13);
			MULT_14(8)<=signed(DIN_14_7)*signed(FMAP_9_14);
			MULT_15(8)<=signed(DIN_15_7)*signed(FMAP_9_15);
			MULT_16(8)<=signed(DIN_16_7)*signed(FMAP_9_16);
			MULT_17(8)<=signed(DIN_17_7)*signed(FMAP_9_17);
			MULT_18(8)<=signed(DIN_18_7)*signed(FMAP_9_18);
			MULT_19(8)<=signed(DIN_19_7)*signed(FMAP_9_19);
			MULT_20(8)<=signed(DIN_20_7)*signed(FMAP_9_20);
			MULT_21(8)<=signed(DIN_21_7)*signed(FMAP_9_21);
			MULT_22(8)<=signed(DIN_22_7)*signed(FMAP_9_22);
			MULT_23(8)<=signed(DIN_23_7)*signed(FMAP_9_23);
			MULT_24(8)<=signed(DIN_24_7)*signed(FMAP_9_24);
			MULT_25(8)<=signed(DIN_25_7)*signed(FMAP_9_25);
			MULT_26(8)<=signed(DIN_26_7)*signed(FMAP_9_26);
			MULT_27(8)<=signed(DIN_27_7)*signed(FMAP_9_27);
			MULT_28(8)<=signed(DIN_28_7)*signed(FMAP_9_28);
			MULT_29(8)<=signed(DIN_29_7)*signed(FMAP_9_29);
			MULT_30(8)<=signed(DIN_30_7)*signed(FMAP_9_30);
			MULT_31(8)<=signed(DIN_31_7)*signed(FMAP_9_31);
			MULT_32(8)<=signed(DIN_32_7)*signed(FMAP_9_32);
			MULT_33(8)<=signed(DIN_33_7)*signed(FMAP_9_33);
			MULT_34(8)<=signed(DIN_34_7)*signed(FMAP_9_34);
			MULT_35(8)<=signed(DIN_35_7)*signed(FMAP_9_35);
			MULT_36(8)<=signed(DIN_36_7)*signed(FMAP_9_36);
			MULT_37(8)<=signed(DIN_37_7)*signed(FMAP_9_37);
			MULT_38(8)<=signed(DIN_38_7)*signed(FMAP_9_38);
			MULT_39(8)<=signed(DIN_39_7)*signed(FMAP_9_39);
			MULT_40(8)<=signed(DIN_40_7)*signed(FMAP_9_40);
			MULT_41(8)<=signed(DIN_41_7)*signed(FMAP_9_41);
			MULT_42(8)<=signed(DIN_42_7)*signed(FMAP_9_42);
			MULT_43(8)<=signed(DIN_43_7)*signed(FMAP_9_43);
			MULT_44(8)<=signed(DIN_44_7)*signed(FMAP_9_44);
			MULT_45(8)<=signed(DIN_45_7)*signed(FMAP_9_45);
			MULT_46(8)<=signed(DIN_46_7)*signed(FMAP_9_46);
			MULT_47(8)<=signed(DIN_47_7)*signed(FMAP_9_47);
			MULT_48(8)<=signed(DIN_48_7)*signed(FMAP_9_48);
			MULT_49(8)<=signed(DIN_49_7)*signed(FMAP_9_49);
			MULT_50(8)<=signed(DIN_50_7)*signed(FMAP_9_50);
			MULT_51(8)<=signed(DIN_51_7)*signed(FMAP_9_51);
			MULT_52(8)<=signed(DIN_52_7)*signed(FMAP_9_52);
			MULT_53(8)<=signed(DIN_53_7)*signed(FMAP_9_53);
			MULT_54(8)<=signed(DIN_54_7)*signed(FMAP_9_54);
			MULT_55(8)<=signed(DIN_55_7)*signed(FMAP_9_55);
			MULT_56(8)<=signed(DIN_56_7)*signed(FMAP_9_56);
			MULT_57(8)<=signed(DIN_57_7)*signed(FMAP_9_57);
			MULT_58(8)<=signed(DIN_58_7)*signed(FMAP_9_58);
			MULT_59(8)<=signed(DIN_59_7)*signed(FMAP_9_59);
			MULT_60(8)<=signed(DIN_60_7)*signed(FMAP_9_60);
			MULT_61(8)<=signed(DIN_61_7)*signed(FMAP_9_61);
			MULT_62(8)<=signed(DIN_62_7)*signed(FMAP_9_62);
			MULT_63(8)<=signed(DIN_63_7)*signed(FMAP_9_63);
			MULT_64(8)<=signed(DIN_64_7)*signed(FMAP_9_64);
			MULT_65(8)<=signed(DIN_65_7)*signed(FMAP_9_65);
			MULT_66(8)<=signed(DIN_66_7)*signed(FMAP_9_66);
			MULT_67(8)<=signed(DIN_67_7)*signed(FMAP_9_67);
			MULT_68(8)<=signed(DIN_68_7)*signed(FMAP_9_68);
			MULT_69(8)<=signed(DIN_69_7)*signed(FMAP_9_69);
			MULT_70(8)<=signed(DIN_70_7)*signed(FMAP_9_70);
			MULT_71(8)<=signed(DIN_71_7)*signed(FMAP_9_71);
			MULT_72(8)<=signed(DIN_72_7)*signed(FMAP_9_72);
			MULT_73(8)<=signed(DIN_73_7)*signed(FMAP_9_73);
			MULT_74(8)<=signed(DIN_74_7)*signed(FMAP_9_74);
			MULT_75(8)<=signed(DIN_75_7)*signed(FMAP_9_75);
			MULT_76(8)<=signed(DIN_76_7)*signed(FMAP_9_76);
			MULT_77(8)<=signed(DIN_77_7)*signed(FMAP_9_77);
			MULT_78(8)<=signed(DIN_78_7)*signed(FMAP_9_78);
			MULT_79(8)<=signed(DIN_79_7)*signed(FMAP_9_79);
			MULT_80(8)<=signed(DIN_80_7)*signed(FMAP_9_80);
			MULT_81(8)<=signed(DIN_81_7)*signed(FMAP_9_81);
			MULT_82(8)<=signed(DIN_82_7)*signed(FMAP_9_82);
			MULT_83(8)<=signed(DIN_83_7)*signed(FMAP_9_83);
			MULT_84(8)<=signed(DIN_84_7)*signed(FMAP_9_84);
			MULT_85(8)<=signed(DIN_85_7)*signed(FMAP_9_85);
			MULT_86(8)<=signed(DIN_86_7)*signed(FMAP_9_86);
			MULT_87(8)<=signed(DIN_87_7)*signed(FMAP_9_87);
			MULT_88(8)<=signed(DIN_88_7)*signed(FMAP_9_88);
			MULT_89(8)<=signed(DIN_89_7)*signed(FMAP_9_89);
			MULT_90(8)<=signed(DIN_90_7)*signed(FMAP_9_90);
			MULT_91(8)<=signed(DIN_91_7)*signed(FMAP_9_91);
			MULT_92(8)<=signed(DIN_92_7)*signed(FMAP_9_92);
			MULT_93(8)<=signed(DIN_93_7)*signed(FMAP_9_93);
			MULT_94(8)<=signed(DIN_94_7)*signed(FMAP_9_94);
			MULT_95(8)<=signed(DIN_95_7)*signed(FMAP_9_95);
			MULT_96(8)<=signed(DIN_96_7)*signed(FMAP_9_96);
			MULT_97(8)<=signed(DIN_97_7)*signed(FMAP_9_97);
			MULT_98(8)<=signed(DIN_98_7)*signed(FMAP_9_98);
			MULT_99(8)<=signed(DIN_99_7)*signed(FMAP_9_99);
			MULT_100(8)<=signed(DIN_100_7)*signed(FMAP_9_100);
			MULT_101(8)<=signed(DIN_101_7)*signed(FMAP_9_101);
			MULT_102(8)<=signed(DIN_102_7)*signed(FMAP_9_102);
			MULT_103(8)<=signed(DIN_103_7)*signed(FMAP_9_103);
			MULT_104(8)<=signed(DIN_104_7)*signed(FMAP_9_104);
			MULT_105(8)<=signed(DIN_105_7)*signed(FMAP_9_105);
			MULT_106(8)<=signed(DIN_106_7)*signed(FMAP_9_106);
			MULT_107(8)<=signed(DIN_107_7)*signed(FMAP_9_107);
			MULT_108(8)<=signed(DIN_108_7)*signed(FMAP_9_108);
			MULT_109(8)<=signed(DIN_109_7)*signed(FMAP_9_109);
			MULT_110(8)<=signed(DIN_110_7)*signed(FMAP_9_110);
			MULT_111(8)<=signed(DIN_111_7)*signed(FMAP_9_111);
			MULT_112(8)<=signed(DIN_112_7)*signed(FMAP_9_112);
			MULT_113(8)<=signed(DIN_113_7)*signed(FMAP_9_113);
			MULT_114(8)<=signed(DIN_114_7)*signed(FMAP_9_114);
			MULT_115(8)<=signed(DIN_115_7)*signed(FMAP_9_115);
			MULT_116(8)<=signed(DIN_116_7)*signed(FMAP_9_116);
			MULT_117(8)<=signed(DIN_117_7)*signed(FMAP_9_117);
			MULT_118(8)<=signed(DIN_118_7)*signed(FMAP_9_118);
			MULT_119(8)<=signed(DIN_119_7)*signed(FMAP_9_119);
			MULT_120(8)<=signed(DIN_120_7)*signed(FMAP_9_120);

			MULT_1(9)<=signed(DIN_1_7)*signed(FMAP_10_1);
			MULT_2(9)<=signed(DIN_2_7)*signed(FMAP_10_2);
			MULT_3(9)<=signed(DIN_3_7)*signed(FMAP_10_3);
			MULT_4(9)<=signed(DIN_4_7)*signed(FMAP_10_4);
			MULT_5(9)<=signed(DIN_5_7)*signed(FMAP_10_5);
			MULT_6(9)<=signed(DIN_6_7)*signed(FMAP_10_6);
			MULT_7(9)<=signed(DIN_7_7)*signed(FMAP_10_7);
			MULT_8(9)<=signed(DIN_8_7)*signed(FMAP_10_8);
			MULT_9(9)<=signed(DIN_9_7)*signed(FMAP_10_9);
			MULT_10(9)<=signed(DIN_10_7)*signed(FMAP_10_10);
			MULT_11(9)<=signed(DIN_11_7)*signed(FMAP_10_11);
			MULT_12(9)<=signed(DIN_12_7)*signed(FMAP_10_12);
			MULT_13(9)<=signed(DIN_13_7)*signed(FMAP_10_13);
			MULT_14(9)<=signed(DIN_14_7)*signed(FMAP_10_14);
			MULT_15(9)<=signed(DIN_15_7)*signed(FMAP_10_15);
			MULT_16(9)<=signed(DIN_16_7)*signed(FMAP_10_16);
			MULT_17(9)<=signed(DIN_17_7)*signed(FMAP_10_17);
			MULT_18(9)<=signed(DIN_18_7)*signed(FMAP_10_18);
			MULT_19(9)<=signed(DIN_19_7)*signed(FMAP_10_19);
			MULT_20(9)<=signed(DIN_20_7)*signed(FMAP_10_20);
			MULT_21(9)<=signed(DIN_21_7)*signed(FMAP_10_21);
			MULT_22(9)<=signed(DIN_22_7)*signed(FMAP_10_22);
			MULT_23(9)<=signed(DIN_23_7)*signed(FMAP_10_23);
			MULT_24(9)<=signed(DIN_24_7)*signed(FMAP_10_24);
			MULT_25(9)<=signed(DIN_25_7)*signed(FMAP_10_25);
			MULT_26(9)<=signed(DIN_26_7)*signed(FMAP_10_26);
			MULT_27(9)<=signed(DIN_27_7)*signed(FMAP_10_27);
			MULT_28(9)<=signed(DIN_28_7)*signed(FMAP_10_28);
			MULT_29(9)<=signed(DIN_29_7)*signed(FMAP_10_29);
			MULT_30(9)<=signed(DIN_30_7)*signed(FMAP_10_30);
			MULT_31(9)<=signed(DIN_31_7)*signed(FMAP_10_31);
			MULT_32(9)<=signed(DIN_32_7)*signed(FMAP_10_32);
			MULT_33(9)<=signed(DIN_33_7)*signed(FMAP_10_33);
			MULT_34(9)<=signed(DIN_34_7)*signed(FMAP_10_34);
			MULT_35(9)<=signed(DIN_35_7)*signed(FMAP_10_35);
			MULT_36(9)<=signed(DIN_36_7)*signed(FMAP_10_36);
			MULT_37(9)<=signed(DIN_37_7)*signed(FMAP_10_37);
			MULT_38(9)<=signed(DIN_38_7)*signed(FMAP_10_38);
			MULT_39(9)<=signed(DIN_39_7)*signed(FMAP_10_39);
			MULT_40(9)<=signed(DIN_40_7)*signed(FMAP_10_40);
			MULT_41(9)<=signed(DIN_41_7)*signed(FMAP_10_41);
			MULT_42(9)<=signed(DIN_42_7)*signed(FMAP_10_42);
			MULT_43(9)<=signed(DIN_43_7)*signed(FMAP_10_43);
			MULT_44(9)<=signed(DIN_44_7)*signed(FMAP_10_44);
			MULT_45(9)<=signed(DIN_45_7)*signed(FMAP_10_45);
			MULT_46(9)<=signed(DIN_46_7)*signed(FMAP_10_46);
			MULT_47(9)<=signed(DIN_47_7)*signed(FMAP_10_47);
			MULT_48(9)<=signed(DIN_48_7)*signed(FMAP_10_48);
			MULT_49(9)<=signed(DIN_49_7)*signed(FMAP_10_49);
			MULT_50(9)<=signed(DIN_50_7)*signed(FMAP_10_50);
			MULT_51(9)<=signed(DIN_51_7)*signed(FMAP_10_51);
			MULT_52(9)<=signed(DIN_52_7)*signed(FMAP_10_52);
			MULT_53(9)<=signed(DIN_53_7)*signed(FMAP_10_53);
			MULT_54(9)<=signed(DIN_54_7)*signed(FMAP_10_54);
			MULT_55(9)<=signed(DIN_55_7)*signed(FMAP_10_55);
			MULT_56(9)<=signed(DIN_56_7)*signed(FMAP_10_56);
			MULT_57(9)<=signed(DIN_57_7)*signed(FMAP_10_57);
			MULT_58(9)<=signed(DIN_58_7)*signed(FMAP_10_58);
			MULT_59(9)<=signed(DIN_59_7)*signed(FMAP_10_59);
			MULT_60(9)<=signed(DIN_60_7)*signed(FMAP_10_60);
			MULT_61(9)<=signed(DIN_61_7)*signed(FMAP_10_61);
			MULT_62(9)<=signed(DIN_62_7)*signed(FMAP_10_62);
			MULT_63(9)<=signed(DIN_63_7)*signed(FMAP_10_63);
			MULT_64(9)<=signed(DIN_64_7)*signed(FMAP_10_64);
			MULT_65(9)<=signed(DIN_65_7)*signed(FMAP_10_65);
			MULT_66(9)<=signed(DIN_66_7)*signed(FMAP_10_66);
			MULT_67(9)<=signed(DIN_67_7)*signed(FMAP_10_67);
			MULT_68(9)<=signed(DIN_68_7)*signed(FMAP_10_68);
			MULT_69(9)<=signed(DIN_69_7)*signed(FMAP_10_69);
			MULT_70(9)<=signed(DIN_70_7)*signed(FMAP_10_70);
			MULT_71(9)<=signed(DIN_71_7)*signed(FMAP_10_71);
			MULT_72(9)<=signed(DIN_72_7)*signed(FMAP_10_72);
			MULT_73(9)<=signed(DIN_73_7)*signed(FMAP_10_73);
			MULT_74(9)<=signed(DIN_74_7)*signed(FMAP_10_74);
			MULT_75(9)<=signed(DIN_75_7)*signed(FMAP_10_75);
			MULT_76(9)<=signed(DIN_76_7)*signed(FMAP_10_76);
			MULT_77(9)<=signed(DIN_77_7)*signed(FMAP_10_77);
			MULT_78(9)<=signed(DIN_78_7)*signed(FMAP_10_78);
			MULT_79(9)<=signed(DIN_79_7)*signed(FMAP_10_79);
			MULT_80(9)<=signed(DIN_80_7)*signed(FMAP_10_80);
			MULT_81(9)<=signed(DIN_81_7)*signed(FMAP_10_81);
			MULT_82(9)<=signed(DIN_82_7)*signed(FMAP_10_82);
			MULT_83(9)<=signed(DIN_83_7)*signed(FMAP_10_83);
			MULT_84(9)<=signed(DIN_84_7)*signed(FMAP_10_84);
			MULT_85(9)<=signed(DIN_85_7)*signed(FMAP_10_85);
			MULT_86(9)<=signed(DIN_86_7)*signed(FMAP_10_86);
			MULT_87(9)<=signed(DIN_87_7)*signed(FMAP_10_87);
			MULT_88(9)<=signed(DIN_88_7)*signed(FMAP_10_88);
			MULT_89(9)<=signed(DIN_89_7)*signed(FMAP_10_89);
			MULT_90(9)<=signed(DIN_90_7)*signed(FMAP_10_90);
			MULT_91(9)<=signed(DIN_91_7)*signed(FMAP_10_91);
			MULT_92(9)<=signed(DIN_92_7)*signed(FMAP_10_92);
			MULT_93(9)<=signed(DIN_93_7)*signed(FMAP_10_93);
			MULT_94(9)<=signed(DIN_94_7)*signed(FMAP_10_94);
			MULT_95(9)<=signed(DIN_95_7)*signed(FMAP_10_95);
			MULT_96(9)<=signed(DIN_96_7)*signed(FMAP_10_96);
			MULT_97(9)<=signed(DIN_97_7)*signed(FMAP_10_97);
			MULT_98(9)<=signed(DIN_98_7)*signed(FMAP_10_98);
			MULT_99(9)<=signed(DIN_99_7)*signed(FMAP_10_99);
			MULT_100(9)<=signed(DIN_100_7)*signed(FMAP_10_100);
			MULT_101(9)<=signed(DIN_101_7)*signed(FMAP_10_101);
			MULT_102(9)<=signed(DIN_102_7)*signed(FMAP_10_102);
			MULT_103(9)<=signed(DIN_103_7)*signed(FMAP_10_103);
			MULT_104(9)<=signed(DIN_104_7)*signed(FMAP_10_104);
			MULT_105(9)<=signed(DIN_105_7)*signed(FMAP_10_105);
			MULT_106(9)<=signed(DIN_106_7)*signed(FMAP_10_106);
			MULT_107(9)<=signed(DIN_107_7)*signed(FMAP_10_107);
			MULT_108(9)<=signed(DIN_108_7)*signed(FMAP_10_108);
			MULT_109(9)<=signed(DIN_109_7)*signed(FMAP_10_109);
			MULT_110(9)<=signed(DIN_110_7)*signed(FMAP_10_110);
			MULT_111(9)<=signed(DIN_111_7)*signed(FMAP_10_111);
			MULT_112(9)<=signed(DIN_112_7)*signed(FMAP_10_112);
			MULT_113(9)<=signed(DIN_113_7)*signed(FMAP_10_113);
			MULT_114(9)<=signed(DIN_114_7)*signed(FMAP_10_114);
			MULT_115(9)<=signed(DIN_115_7)*signed(FMAP_10_115);
			MULT_116(9)<=signed(DIN_116_7)*signed(FMAP_10_116);
			MULT_117(9)<=signed(DIN_117_7)*signed(FMAP_10_117);
			MULT_118(9)<=signed(DIN_118_7)*signed(FMAP_10_118);
			MULT_119(9)<=signed(DIN_119_7)*signed(FMAP_10_119);
			MULT_120(9)<=signed(DIN_120_7)*signed(FMAP_10_120);

			MULT_1(10)<=signed(DIN_1_7)*signed(FMAP_11_1);
			MULT_2(10)<=signed(DIN_2_7)*signed(FMAP_11_2);
			MULT_3(10)<=signed(DIN_3_7)*signed(FMAP_11_3);
			MULT_4(10)<=signed(DIN_4_7)*signed(FMAP_11_4);
			MULT_5(10)<=signed(DIN_5_7)*signed(FMAP_11_5);
			MULT_6(10)<=signed(DIN_6_7)*signed(FMAP_11_6);
			MULT_7(10)<=signed(DIN_7_7)*signed(FMAP_11_7);
			MULT_8(10)<=signed(DIN_8_7)*signed(FMAP_11_8);
			MULT_9(10)<=signed(DIN_9_7)*signed(FMAP_11_9);
			MULT_10(10)<=signed(DIN_10_7)*signed(FMAP_11_10);
			MULT_11(10)<=signed(DIN_11_7)*signed(FMAP_11_11);
			MULT_12(10)<=signed(DIN_12_7)*signed(FMAP_11_12);
			MULT_13(10)<=signed(DIN_13_7)*signed(FMAP_11_13);
			MULT_14(10)<=signed(DIN_14_7)*signed(FMAP_11_14);
			MULT_15(10)<=signed(DIN_15_7)*signed(FMAP_11_15);
			MULT_16(10)<=signed(DIN_16_7)*signed(FMAP_11_16);
			MULT_17(10)<=signed(DIN_17_7)*signed(FMAP_11_17);
			MULT_18(10)<=signed(DIN_18_7)*signed(FMAP_11_18);
			MULT_19(10)<=signed(DIN_19_7)*signed(FMAP_11_19);
			MULT_20(10)<=signed(DIN_20_7)*signed(FMAP_11_20);
			MULT_21(10)<=signed(DIN_21_7)*signed(FMAP_11_21);
			MULT_22(10)<=signed(DIN_22_7)*signed(FMAP_11_22);
			MULT_23(10)<=signed(DIN_23_7)*signed(FMAP_11_23);
			MULT_24(10)<=signed(DIN_24_7)*signed(FMAP_11_24);
			MULT_25(10)<=signed(DIN_25_7)*signed(FMAP_11_25);
			MULT_26(10)<=signed(DIN_26_7)*signed(FMAP_11_26);
			MULT_27(10)<=signed(DIN_27_7)*signed(FMAP_11_27);
			MULT_28(10)<=signed(DIN_28_7)*signed(FMAP_11_28);
			MULT_29(10)<=signed(DIN_29_7)*signed(FMAP_11_29);
			MULT_30(10)<=signed(DIN_30_7)*signed(FMAP_11_30);
			MULT_31(10)<=signed(DIN_31_7)*signed(FMAP_11_31);
			MULT_32(10)<=signed(DIN_32_7)*signed(FMAP_11_32);
			MULT_33(10)<=signed(DIN_33_7)*signed(FMAP_11_33);
			MULT_34(10)<=signed(DIN_34_7)*signed(FMAP_11_34);
			MULT_35(10)<=signed(DIN_35_7)*signed(FMAP_11_35);
			MULT_36(10)<=signed(DIN_36_7)*signed(FMAP_11_36);
			MULT_37(10)<=signed(DIN_37_7)*signed(FMAP_11_37);
			MULT_38(10)<=signed(DIN_38_7)*signed(FMAP_11_38);
			MULT_39(10)<=signed(DIN_39_7)*signed(FMAP_11_39);
			MULT_40(10)<=signed(DIN_40_7)*signed(FMAP_11_40);
			MULT_41(10)<=signed(DIN_41_7)*signed(FMAP_11_41);
			MULT_42(10)<=signed(DIN_42_7)*signed(FMAP_11_42);
			MULT_43(10)<=signed(DIN_43_7)*signed(FMAP_11_43);
			MULT_44(10)<=signed(DIN_44_7)*signed(FMAP_11_44);
			MULT_45(10)<=signed(DIN_45_7)*signed(FMAP_11_45);
			MULT_46(10)<=signed(DIN_46_7)*signed(FMAP_11_46);
			MULT_47(10)<=signed(DIN_47_7)*signed(FMAP_11_47);
			MULT_48(10)<=signed(DIN_48_7)*signed(FMAP_11_48);
			MULT_49(10)<=signed(DIN_49_7)*signed(FMAP_11_49);
			MULT_50(10)<=signed(DIN_50_7)*signed(FMAP_11_50);
			MULT_51(10)<=signed(DIN_51_7)*signed(FMAP_11_51);
			MULT_52(10)<=signed(DIN_52_7)*signed(FMAP_11_52);
			MULT_53(10)<=signed(DIN_53_7)*signed(FMAP_11_53);
			MULT_54(10)<=signed(DIN_54_7)*signed(FMAP_11_54);
			MULT_55(10)<=signed(DIN_55_7)*signed(FMAP_11_55);
			MULT_56(10)<=signed(DIN_56_7)*signed(FMAP_11_56);
			MULT_57(10)<=signed(DIN_57_7)*signed(FMAP_11_57);
			MULT_58(10)<=signed(DIN_58_7)*signed(FMAP_11_58);
			MULT_59(10)<=signed(DIN_59_7)*signed(FMAP_11_59);
			MULT_60(10)<=signed(DIN_60_7)*signed(FMAP_11_60);
			MULT_61(10)<=signed(DIN_61_7)*signed(FMAP_11_61);
			MULT_62(10)<=signed(DIN_62_7)*signed(FMAP_11_62);
			MULT_63(10)<=signed(DIN_63_7)*signed(FMAP_11_63);
			MULT_64(10)<=signed(DIN_64_7)*signed(FMAP_11_64);
			MULT_65(10)<=signed(DIN_65_7)*signed(FMAP_11_65);
			MULT_66(10)<=signed(DIN_66_7)*signed(FMAP_11_66);
			MULT_67(10)<=signed(DIN_67_7)*signed(FMAP_11_67);
			MULT_68(10)<=signed(DIN_68_7)*signed(FMAP_11_68);
			MULT_69(10)<=signed(DIN_69_7)*signed(FMAP_11_69);
			MULT_70(10)<=signed(DIN_70_7)*signed(FMAP_11_70);
			MULT_71(10)<=signed(DIN_71_7)*signed(FMAP_11_71);
			MULT_72(10)<=signed(DIN_72_7)*signed(FMAP_11_72);
			MULT_73(10)<=signed(DIN_73_7)*signed(FMAP_11_73);
			MULT_74(10)<=signed(DIN_74_7)*signed(FMAP_11_74);
			MULT_75(10)<=signed(DIN_75_7)*signed(FMAP_11_75);
			MULT_76(10)<=signed(DIN_76_7)*signed(FMAP_11_76);
			MULT_77(10)<=signed(DIN_77_7)*signed(FMAP_11_77);
			MULT_78(10)<=signed(DIN_78_7)*signed(FMAP_11_78);
			MULT_79(10)<=signed(DIN_79_7)*signed(FMAP_11_79);
			MULT_80(10)<=signed(DIN_80_7)*signed(FMAP_11_80);
			MULT_81(10)<=signed(DIN_81_7)*signed(FMAP_11_81);
			MULT_82(10)<=signed(DIN_82_7)*signed(FMAP_11_82);
			MULT_83(10)<=signed(DIN_83_7)*signed(FMAP_11_83);
			MULT_84(10)<=signed(DIN_84_7)*signed(FMAP_11_84);
			MULT_85(10)<=signed(DIN_85_7)*signed(FMAP_11_85);
			MULT_86(10)<=signed(DIN_86_7)*signed(FMAP_11_86);
			MULT_87(10)<=signed(DIN_87_7)*signed(FMAP_11_87);
			MULT_88(10)<=signed(DIN_88_7)*signed(FMAP_11_88);
			MULT_89(10)<=signed(DIN_89_7)*signed(FMAP_11_89);
			MULT_90(10)<=signed(DIN_90_7)*signed(FMAP_11_90);
			MULT_91(10)<=signed(DIN_91_7)*signed(FMAP_11_91);
			MULT_92(10)<=signed(DIN_92_7)*signed(FMAP_11_92);
			MULT_93(10)<=signed(DIN_93_7)*signed(FMAP_11_93);
			MULT_94(10)<=signed(DIN_94_7)*signed(FMAP_11_94);
			MULT_95(10)<=signed(DIN_95_7)*signed(FMAP_11_95);
			MULT_96(10)<=signed(DIN_96_7)*signed(FMAP_11_96);
			MULT_97(10)<=signed(DIN_97_7)*signed(FMAP_11_97);
			MULT_98(10)<=signed(DIN_98_7)*signed(FMAP_11_98);
			MULT_99(10)<=signed(DIN_99_7)*signed(FMAP_11_99);
			MULT_100(10)<=signed(DIN_100_7)*signed(FMAP_11_100);
			MULT_101(10)<=signed(DIN_101_7)*signed(FMAP_11_101);
			MULT_102(10)<=signed(DIN_102_7)*signed(FMAP_11_102);
			MULT_103(10)<=signed(DIN_103_7)*signed(FMAP_11_103);
			MULT_104(10)<=signed(DIN_104_7)*signed(FMAP_11_104);
			MULT_105(10)<=signed(DIN_105_7)*signed(FMAP_11_105);
			MULT_106(10)<=signed(DIN_106_7)*signed(FMAP_11_106);
			MULT_107(10)<=signed(DIN_107_7)*signed(FMAP_11_107);
			MULT_108(10)<=signed(DIN_108_7)*signed(FMAP_11_108);
			MULT_109(10)<=signed(DIN_109_7)*signed(FMAP_11_109);
			MULT_110(10)<=signed(DIN_110_7)*signed(FMAP_11_110);
			MULT_111(10)<=signed(DIN_111_7)*signed(FMAP_11_111);
			MULT_112(10)<=signed(DIN_112_7)*signed(FMAP_11_112);
			MULT_113(10)<=signed(DIN_113_7)*signed(FMAP_11_113);
			MULT_114(10)<=signed(DIN_114_7)*signed(FMAP_11_114);
			MULT_115(10)<=signed(DIN_115_7)*signed(FMAP_11_115);
			MULT_116(10)<=signed(DIN_116_7)*signed(FMAP_11_116);
			MULT_117(10)<=signed(DIN_117_7)*signed(FMAP_11_117);
			MULT_118(10)<=signed(DIN_118_7)*signed(FMAP_11_118);
			MULT_119(10)<=signed(DIN_119_7)*signed(FMAP_11_119);
			MULT_120(10)<=signed(DIN_120_7)*signed(FMAP_11_120);

			MULT_1(11)<=signed(DIN_1_7)*signed(FMAP_12_1);
			MULT_2(11)<=signed(DIN_2_7)*signed(FMAP_12_2);
			MULT_3(11)<=signed(DIN_3_7)*signed(FMAP_12_3);
			MULT_4(11)<=signed(DIN_4_7)*signed(FMAP_12_4);
			MULT_5(11)<=signed(DIN_5_7)*signed(FMAP_12_5);
			MULT_6(11)<=signed(DIN_6_7)*signed(FMAP_12_6);
			MULT_7(11)<=signed(DIN_7_7)*signed(FMAP_12_7);
			MULT_8(11)<=signed(DIN_8_7)*signed(FMAP_12_8);
			MULT_9(11)<=signed(DIN_9_7)*signed(FMAP_12_9);
			MULT_10(11)<=signed(DIN_10_7)*signed(FMAP_12_10);
			MULT_11(11)<=signed(DIN_11_7)*signed(FMAP_12_11);
			MULT_12(11)<=signed(DIN_12_7)*signed(FMAP_12_12);
			MULT_13(11)<=signed(DIN_13_7)*signed(FMAP_12_13);
			MULT_14(11)<=signed(DIN_14_7)*signed(FMAP_12_14);
			MULT_15(11)<=signed(DIN_15_7)*signed(FMAP_12_15);
			MULT_16(11)<=signed(DIN_16_7)*signed(FMAP_12_16);
			MULT_17(11)<=signed(DIN_17_7)*signed(FMAP_12_17);
			MULT_18(11)<=signed(DIN_18_7)*signed(FMAP_12_18);
			MULT_19(11)<=signed(DIN_19_7)*signed(FMAP_12_19);
			MULT_20(11)<=signed(DIN_20_7)*signed(FMAP_12_20);
			MULT_21(11)<=signed(DIN_21_7)*signed(FMAP_12_21);
			MULT_22(11)<=signed(DIN_22_7)*signed(FMAP_12_22);
			MULT_23(11)<=signed(DIN_23_7)*signed(FMAP_12_23);
			MULT_24(11)<=signed(DIN_24_7)*signed(FMAP_12_24);
			MULT_25(11)<=signed(DIN_25_7)*signed(FMAP_12_25);
			MULT_26(11)<=signed(DIN_26_7)*signed(FMAP_12_26);
			MULT_27(11)<=signed(DIN_27_7)*signed(FMAP_12_27);
			MULT_28(11)<=signed(DIN_28_7)*signed(FMAP_12_28);
			MULT_29(11)<=signed(DIN_29_7)*signed(FMAP_12_29);
			MULT_30(11)<=signed(DIN_30_7)*signed(FMAP_12_30);
			MULT_31(11)<=signed(DIN_31_7)*signed(FMAP_12_31);
			MULT_32(11)<=signed(DIN_32_7)*signed(FMAP_12_32);
			MULT_33(11)<=signed(DIN_33_7)*signed(FMAP_12_33);
			MULT_34(11)<=signed(DIN_34_7)*signed(FMAP_12_34);
			MULT_35(11)<=signed(DIN_35_7)*signed(FMAP_12_35);
			MULT_36(11)<=signed(DIN_36_7)*signed(FMAP_12_36);
			MULT_37(11)<=signed(DIN_37_7)*signed(FMAP_12_37);
			MULT_38(11)<=signed(DIN_38_7)*signed(FMAP_12_38);
			MULT_39(11)<=signed(DIN_39_7)*signed(FMAP_12_39);
			MULT_40(11)<=signed(DIN_40_7)*signed(FMAP_12_40);
			MULT_41(11)<=signed(DIN_41_7)*signed(FMAP_12_41);
			MULT_42(11)<=signed(DIN_42_7)*signed(FMAP_12_42);
			MULT_43(11)<=signed(DIN_43_7)*signed(FMAP_12_43);
			MULT_44(11)<=signed(DIN_44_7)*signed(FMAP_12_44);
			MULT_45(11)<=signed(DIN_45_7)*signed(FMAP_12_45);
			MULT_46(11)<=signed(DIN_46_7)*signed(FMAP_12_46);
			MULT_47(11)<=signed(DIN_47_7)*signed(FMAP_12_47);
			MULT_48(11)<=signed(DIN_48_7)*signed(FMAP_12_48);
			MULT_49(11)<=signed(DIN_49_7)*signed(FMAP_12_49);
			MULT_50(11)<=signed(DIN_50_7)*signed(FMAP_12_50);
			MULT_51(11)<=signed(DIN_51_7)*signed(FMAP_12_51);
			MULT_52(11)<=signed(DIN_52_7)*signed(FMAP_12_52);
			MULT_53(11)<=signed(DIN_53_7)*signed(FMAP_12_53);
			MULT_54(11)<=signed(DIN_54_7)*signed(FMAP_12_54);
			MULT_55(11)<=signed(DIN_55_7)*signed(FMAP_12_55);
			MULT_56(11)<=signed(DIN_56_7)*signed(FMAP_12_56);
			MULT_57(11)<=signed(DIN_57_7)*signed(FMAP_12_57);
			MULT_58(11)<=signed(DIN_58_7)*signed(FMAP_12_58);
			MULT_59(11)<=signed(DIN_59_7)*signed(FMAP_12_59);
			MULT_60(11)<=signed(DIN_60_7)*signed(FMAP_12_60);
			MULT_61(11)<=signed(DIN_61_7)*signed(FMAP_12_61);
			MULT_62(11)<=signed(DIN_62_7)*signed(FMAP_12_62);
			MULT_63(11)<=signed(DIN_63_7)*signed(FMAP_12_63);
			MULT_64(11)<=signed(DIN_64_7)*signed(FMAP_12_64);
			MULT_65(11)<=signed(DIN_65_7)*signed(FMAP_12_65);
			MULT_66(11)<=signed(DIN_66_7)*signed(FMAP_12_66);
			MULT_67(11)<=signed(DIN_67_7)*signed(FMAP_12_67);
			MULT_68(11)<=signed(DIN_68_7)*signed(FMAP_12_68);
			MULT_69(11)<=signed(DIN_69_7)*signed(FMAP_12_69);
			MULT_70(11)<=signed(DIN_70_7)*signed(FMAP_12_70);
			MULT_71(11)<=signed(DIN_71_7)*signed(FMAP_12_71);
			MULT_72(11)<=signed(DIN_72_7)*signed(FMAP_12_72);
			MULT_73(11)<=signed(DIN_73_7)*signed(FMAP_12_73);
			MULT_74(11)<=signed(DIN_74_7)*signed(FMAP_12_74);
			MULT_75(11)<=signed(DIN_75_7)*signed(FMAP_12_75);
			MULT_76(11)<=signed(DIN_76_7)*signed(FMAP_12_76);
			MULT_77(11)<=signed(DIN_77_7)*signed(FMAP_12_77);
			MULT_78(11)<=signed(DIN_78_7)*signed(FMAP_12_78);
			MULT_79(11)<=signed(DIN_79_7)*signed(FMAP_12_79);
			MULT_80(11)<=signed(DIN_80_7)*signed(FMAP_12_80);
			MULT_81(11)<=signed(DIN_81_7)*signed(FMAP_12_81);
			MULT_82(11)<=signed(DIN_82_7)*signed(FMAP_12_82);
			MULT_83(11)<=signed(DIN_83_7)*signed(FMAP_12_83);
			MULT_84(11)<=signed(DIN_84_7)*signed(FMAP_12_84);
			MULT_85(11)<=signed(DIN_85_7)*signed(FMAP_12_85);
			MULT_86(11)<=signed(DIN_86_7)*signed(FMAP_12_86);
			MULT_87(11)<=signed(DIN_87_7)*signed(FMAP_12_87);
			MULT_88(11)<=signed(DIN_88_7)*signed(FMAP_12_88);
			MULT_89(11)<=signed(DIN_89_7)*signed(FMAP_12_89);
			MULT_90(11)<=signed(DIN_90_7)*signed(FMAP_12_90);
			MULT_91(11)<=signed(DIN_91_7)*signed(FMAP_12_91);
			MULT_92(11)<=signed(DIN_92_7)*signed(FMAP_12_92);
			MULT_93(11)<=signed(DIN_93_7)*signed(FMAP_12_93);
			MULT_94(11)<=signed(DIN_94_7)*signed(FMAP_12_94);
			MULT_95(11)<=signed(DIN_95_7)*signed(FMAP_12_95);
			MULT_96(11)<=signed(DIN_96_7)*signed(FMAP_12_96);
			MULT_97(11)<=signed(DIN_97_7)*signed(FMAP_12_97);
			MULT_98(11)<=signed(DIN_98_7)*signed(FMAP_12_98);
			MULT_99(11)<=signed(DIN_99_7)*signed(FMAP_12_99);
			MULT_100(11)<=signed(DIN_100_7)*signed(FMAP_12_100);
			MULT_101(11)<=signed(DIN_101_7)*signed(FMAP_12_101);
			MULT_102(11)<=signed(DIN_102_7)*signed(FMAP_12_102);
			MULT_103(11)<=signed(DIN_103_7)*signed(FMAP_12_103);
			MULT_104(11)<=signed(DIN_104_7)*signed(FMAP_12_104);
			MULT_105(11)<=signed(DIN_105_7)*signed(FMAP_12_105);
			MULT_106(11)<=signed(DIN_106_7)*signed(FMAP_12_106);
			MULT_107(11)<=signed(DIN_107_7)*signed(FMAP_12_107);
			MULT_108(11)<=signed(DIN_108_7)*signed(FMAP_12_108);
			MULT_109(11)<=signed(DIN_109_7)*signed(FMAP_12_109);
			MULT_110(11)<=signed(DIN_110_7)*signed(FMAP_12_110);
			MULT_111(11)<=signed(DIN_111_7)*signed(FMAP_12_111);
			MULT_112(11)<=signed(DIN_112_7)*signed(FMAP_12_112);
			MULT_113(11)<=signed(DIN_113_7)*signed(FMAP_12_113);
			MULT_114(11)<=signed(DIN_114_7)*signed(FMAP_12_114);
			MULT_115(11)<=signed(DIN_115_7)*signed(FMAP_12_115);
			MULT_116(11)<=signed(DIN_116_7)*signed(FMAP_12_116);
			MULT_117(11)<=signed(DIN_117_7)*signed(FMAP_12_117);
			MULT_118(11)<=signed(DIN_118_7)*signed(FMAP_12_118);
			MULT_119(11)<=signed(DIN_119_7)*signed(FMAP_12_119);
			MULT_120(11)<=signed(DIN_120_7)*signed(FMAP_12_120);

			MULT_1(12)<=signed(DIN_1_7)*signed(FMAP_13_1);
			MULT_2(12)<=signed(DIN_2_7)*signed(FMAP_13_2);
			MULT_3(12)<=signed(DIN_3_7)*signed(FMAP_13_3);
			MULT_4(12)<=signed(DIN_4_7)*signed(FMAP_13_4);
			MULT_5(12)<=signed(DIN_5_7)*signed(FMAP_13_5);
			MULT_6(12)<=signed(DIN_6_7)*signed(FMAP_13_6);
			MULT_7(12)<=signed(DIN_7_7)*signed(FMAP_13_7);
			MULT_8(12)<=signed(DIN_8_7)*signed(FMAP_13_8);
			MULT_9(12)<=signed(DIN_9_7)*signed(FMAP_13_9);
			MULT_10(12)<=signed(DIN_10_7)*signed(FMAP_13_10);
			MULT_11(12)<=signed(DIN_11_7)*signed(FMAP_13_11);
			MULT_12(12)<=signed(DIN_12_7)*signed(FMAP_13_12);
			MULT_13(12)<=signed(DIN_13_7)*signed(FMAP_13_13);
			MULT_14(12)<=signed(DIN_14_7)*signed(FMAP_13_14);
			MULT_15(12)<=signed(DIN_15_7)*signed(FMAP_13_15);
			MULT_16(12)<=signed(DIN_16_7)*signed(FMAP_13_16);
			MULT_17(12)<=signed(DIN_17_7)*signed(FMAP_13_17);
			MULT_18(12)<=signed(DIN_18_7)*signed(FMAP_13_18);
			MULT_19(12)<=signed(DIN_19_7)*signed(FMAP_13_19);
			MULT_20(12)<=signed(DIN_20_7)*signed(FMAP_13_20);
			MULT_21(12)<=signed(DIN_21_7)*signed(FMAP_13_21);
			MULT_22(12)<=signed(DIN_22_7)*signed(FMAP_13_22);
			MULT_23(12)<=signed(DIN_23_7)*signed(FMAP_13_23);
			MULT_24(12)<=signed(DIN_24_7)*signed(FMAP_13_24);
			MULT_25(12)<=signed(DIN_25_7)*signed(FMAP_13_25);
			MULT_26(12)<=signed(DIN_26_7)*signed(FMAP_13_26);
			MULT_27(12)<=signed(DIN_27_7)*signed(FMAP_13_27);
			MULT_28(12)<=signed(DIN_28_7)*signed(FMAP_13_28);
			MULT_29(12)<=signed(DIN_29_7)*signed(FMAP_13_29);
			MULT_30(12)<=signed(DIN_30_7)*signed(FMAP_13_30);
			MULT_31(12)<=signed(DIN_31_7)*signed(FMAP_13_31);
			MULT_32(12)<=signed(DIN_32_7)*signed(FMAP_13_32);
			MULT_33(12)<=signed(DIN_33_7)*signed(FMAP_13_33);
			MULT_34(12)<=signed(DIN_34_7)*signed(FMAP_13_34);
			MULT_35(12)<=signed(DIN_35_7)*signed(FMAP_13_35);
			MULT_36(12)<=signed(DIN_36_7)*signed(FMAP_13_36);
			MULT_37(12)<=signed(DIN_37_7)*signed(FMAP_13_37);
			MULT_38(12)<=signed(DIN_38_7)*signed(FMAP_13_38);
			MULT_39(12)<=signed(DIN_39_7)*signed(FMAP_13_39);
			MULT_40(12)<=signed(DIN_40_7)*signed(FMAP_13_40);
			MULT_41(12)<=signed(DIN_41_7)*signed(FMAP_13_41);
			MULT_42(12)<=signed(DIN_42_7)*signed(FMAP_13_42);
			MULT_43(12)<=signed(DIN_43_7)*signed(FMAP_13_43);
			MULT_44(12)<=signed(DIN_44_7)*signed(FMAP_13_44);
			MULT_45(12)<=signed(DIN_45_7)*signed(FMAP_13_45);
			MULT_46(12)<=signed(DIN_46_7)*signed(FMAP_13_46);
			MULT_47(12)<=signed(DIN_47_7)*signed(FMAP_13_47);
			MULT_48(12)<=signed(DIN_48_7)*signed(FMAP_13_48);
			MULT_49(12)<=signed(DIN_49_7)*signed(FMAP_13_49);
			MULT_50(12)<=signed(DIN_50_7)*signed(FMAP_13_50);
			MULT_51(12)<=signed(DIN_51_7)*signed(FMAP_13_51);
			MULT_52(12)<=signed(DIN_52_7)*signed(FMAP_13_52);
			MULT_53(12)<=signed(DIN_53_7)*signed(FMAP_13_53);
			MULT_54(12)<=signed(DIN_54_7)*signed(FMAP_13_54);
			MULT_55(12)<=signed(DIN_55_7)*signed(FMAP_13_55);
			MULT_56(12)<=signed(DIN_56_7)*signed(FMAP_13_56);
			MULT_57(12)<=signed(DIN_57_7)*signed(FMAP_13_57);
			MULT_58(12)<=signed(DIN_58_7)*signed(FMAP_13_58);
			MULT_59(12)<=signed(DIN_59_7)*signed(FMAP_13_59);
			MULT_60(12)<=signed(DIN_60_7)*signed(FMAP_13_60);
			MULT_61(12)<=signed(DIN_61_7)*signed(FMAP_13_61);
			MULT_62(12)<=signed(DIN_62_7)*signed(FMAP_13_62);
			MULT_63(12)<=signed(DIN_63_7)*signed(FMAP_13_63);
			MULT_64(12)<=signed(DIN_64_7)*signed(FMAP_13_64);
			MULT_65(12)<=signed(DIN_65_7)*signed(FMAP_13_65);
			MULT_66(12)<=signed(DIN_66_7)*signed(FMAP_13_66);
			MULT_67(12)<=signed(DIN_67_7)*signed(FMAP_13_67);
			MULT_68(12)<=signed(DIN_68_7)*signed(FMAP_13_68);
			MULT_69(12)<=signed(DIN_69_7)*signed(FMAP_13_69);
			MULT_70(12)<=signed(DIN_70_7)*signed(FMAP_13_70);
			MULT_71(12)<=signed(DIN_71_7)*signed(FMAP_13_71);
			MULT_72(12)<=signed(DIN_72_7)*signed(FMAP_13_72);
			MULT_73(12)<=signed(DIN_73_7)*signed(FMAP_13_73);
			MULT_74(12)<=signed(DIN_74_7)*signed(FMAP_13_74);
			MULT_75(12)<=signed(DIN_75_7)*signed(FMAP_13_75);
			MULT_76(12)<=signed(DIN_76_7)*signed(FMAP_13_76);
			MULT_77(12)<=signed(DIN_77_7)*signed(FMAP_13_77);
			MULT_78(12)<=signed(DIN_78_7)*signed(FMAP_13_78);
			MULT_79(12)<=signed(DIN_79_7)*signed(FMAP_13_79);
			MULT_80(12)<=signed(DIN_80_7)*signed(FMAP_13_80);
			MULT_81(12)<=signed(DIN_81_7)*signed(FMAP_13_81);
			MULT_82(12)<=signed(DIN_82_7)*signed(FMAP_13_82);
			MULT_83(12)<=signed(DIN_83_7)*signed(FMAP_13_83);
			MULT_84(12)<=signed(DIN_84_7)*signed(FMAP_13_84);
			MULT_85(12)<=signed(DIN_85_7)*signed(FMAP_13_85);
			MULT_86(12)<=signed(DIN_86_7)*signed(FMAP_13_86);
			MULT_87(12)<=signed(DIN_87_7)*signed(FMAP_13_87);
			MULT_88(12)<=signed(DIN_88_7)*signed(FMAP_13_88);
			MULT_89(12)<=signed(DIN_89_7)*signed(FMAP_13_89);
			MULT_90(12)<=signed(DIN_90_7)*signed(FMAP_13_90);
			MULT_91(12)<=signed(DIN_91_7)*signed(FMAP_13_91);
			MULT_92(12)<=signed(DIN_92_7)*signed(FMAP_13_92);
			MULT_93(12)<=signed(DIN_93_7)*signed(FMAP_13_93);
			MULT_94(12)<=signed(DIN_94_7)*signed(FMAP_13_94);
			MULT_95(12)<=signed(DIN_95_7)*signed(FMAP_13_95);
			MULT_96(12)<=signed(DIN_96_7)*signed(FMAP_13_96);
			MULT_97(12)<=signed(DIN_97_7)*signed(FMAP_13_97);
			MULT_98(12)<=signed(DIN_98_7)*signed(FMAP_13_98);
			MULT_99(12)<=signed(DIN_99_7)*signed(FMAP_13_99);
			MULT_100(12)<=signed(DIN_100_7)*signed(FMAP_13_100);
			MULT_101(12)<=signed(DIN_101_7)*signed(FMAP_13_101);
			MULT_102(12)<=signed(DIN_102_7)*signed(FMAP_13_102);
			MULT_103(12)<=signed(DIN_103_7)*signed(FMAP_13_103);
			MULT_104(12)<=signed(DIN_104_7)*signed(FMAP_13_104);
			MULT_105(12)<=signed(DIN_105_7)*signed(FMAP_13_105);
			MULT_106(12)<=signed(DIN_106_7)*signed(FMAP_13_106);
			MULT_107(12)<=signed(DIN_107_7)*signed(FMAP_13_107);
			MULT_108(12)<=signed(DIN_108_7)*signed(FMAP_13_108);
			MULT_109(12)<=signed(DIN_109_7)*signed(FMAP_13_109);
			MULT_110(12)<=signed(DIN_110_7)*signed(FMAP_13_110);
			MULT_111(12)<=signed(DIN_111_7)*signed(FMAP_13_111);
			MULT_112(12)<=signed(DIN_112_7)*signed(FMAP_13_112);
			MULT_113(12)<=signed(DIN_113_7)*signed(FMAP_13_113);
			MULT_114(12)<=signed(DIN_114_7)*signed(FMAP_13_114);
			MULT_115(12)<=signed(DIN_115_7)*signed(FMAP_13_115);
			MULT_116(12)<=signed(DIN_116_7)*signed(FMAP_13_116);
			MULT_117(12)<=signed(DIN_117_7)*signed(FMAP_13_117);
			MULT_118(12)<=signed(DIN_118_7)*signed(FMAP_13_118);
			MULT_119(12)<=signed(DIN_119_7)*signed(FMAP_13_119);
			MULT_120(12)<=signed(DIN_120_7)*signed(FMAP_13_120);

			MULT_1(13)<=signed(DIN_1_7)*signed(FMAP_14_1);
			MULT_2(13)<=signed(DIN_2_7)*signed(FMAP_14_2);
			MULT_3(13)<=signed(DIN_3_7)*signed(FMAP_14_3);
			MULT_4(13)<=signed(DIN_4_7)*signed(FMAP_14_4);
			MULT_5(13)<=signed(DIN_5_7)*signed(FMAP_14_5);
			MULT_6(13)<=signed(DIN_6_7)*signed(FMAP_14_6);
			MULT_7(13)<=signed(DIN_7_7)*signed(FMAP_14_7);
			MULT_8(13)<=signed(DIN_8_7)*signed(FMAP_14_8);
			MULT_9(13)<=signed(DIN_9_7)*signed(FMAP_14_9);
			MULT_10(13)<=signed(DIN_10_7)*signed(FMAP_14_10);
			MULT_11(13)<=signed(DIN_11_7)*signed(FMAP_14_11);
			MULT_12(13)<=signed(DIN_12_7)*signed(FMAP_14_12);
			MULT_13(13)<=signed(DIN_13_7)*signed(FMAP_14_13);
			MULT_14(13)<=signed(DIN_14_7)*signed(FMAP_14_14);
			MULT_15(13)<=signed(DIN_15_7)*signed(FMAP_14_15);
			MULT_16(13)<=signed(DIN_16_7)*signed(FMAP_14_16);
			MULT_17(13)<=signed(DIN_17_7)*signed(FMAP_14_17);
			MULT_18(13)<=signed(DIN_18_7)*signed(FMAP_14_18);
			MULT_19(13)<=signed(DIN_19_7)*signed(FMAP_14_19);
			MULT_20(13)<=signed(DIN_20_7)*signed(FMAP_14_20);
			MULT_21(13)<=signed(DIN_21_7)*signed(FMAP_14_21);
			MULT_22(13)<=signed(DIN_22_7)*signed(FMAP_14_22);
			MULT_23(13)<=signed(DIN_23_7)*signed(FMAP_14_23);
			MULT_24(13)<=signed(DIN_24_7)*signed(FMAP_14_24);
			MULT_25(13)<=signed(DIN_25_7)*signed(FMAP_14_25);
			MULT_26(13)<=signed(DIN_26_7)*signed(FMAP_14_26);
			MULT_27(13)<=signed(DIN_27_7)*signed(FMAP_14_27);
			MULT_28(13)<=signed(DIN_28_7)*signed(FMAP_14_28);
			MULT_29(13)<=signed(DIN_29_7)*signed(FMAP_14_29);
			MULT_30(13)<=signed(DIN_30_7)*signed(FMAP_14_30);
			MULT_31(13)<=signed(DIN_31_7)*signed(FMAP_14_31);
			MULT_32(13)<=signed(DIN_32_7)*signed(FMAP_14_32);
			MULT_33(13)<=signed(DIN_33_7)*signed(FMAP_14_33);
			MULT_34(13)<=signed(DIN_34_7)*signed(FMAP_14_34);
			MULT_35(13)<=signed(DIN_35_7)*signed(FMAP_14_35);
			MULT_36(13)<=signed(DIN_36_7)*signed(FMAP_14_36);
			MULT_37(13)<=signed(DIN_37_7)*signed(FMAP_14_37);
			MULT_38(13)<=signed(DIN_38_7)*signed(FMAP_14_38);
			MULT_39(13)<=signed(DIN_39_7)*signed(FMAP_14_39);
			MULT_40(13)<=signed(DIN_40_7)*signed(FMAP_14_40);
			MULT_41(13)<=signed(DIN_41_7)*signed(FMAP_14_41);
			MULT_42(13)<=signed(DIN_42_7)*signed(FMAP_14_42);
			MULT_43(13)<=signed(DIN_43_7)*signed(FMAP_14_43);
			MULT_44(13)<=signed(DIN_44_7)*signed(FMAP_14_44);
			MULT_45(13)<=signed(DIN_45_7)*signed(FMAP_14_45);
			MULT_46(13)<=signed(DIN_46_7)*signed(FMAP_14_46);
			MULT_47(13)<=signed(DIN_47_7)*signed(FMAP_14_47);
			MULT_48(13)<=signed(DIN_48_7)*signed(FMAP_14_48);
			MULT_49(13)<=signed(DIN_49_7)*signed(FMAP_14_49);
			MULT_50(13)<=signed(DIN_50_7)*signed(FMAP_14_50);
			MULT_51(13)<=signed(DIN_51_7)*signed(FMAP_14_51);
			MULT_52(13)<=signed(DIN_52_7)*signed(FMAP_14_52);
			MULT_53(13)<=signed(DIN_53_7)*signed(FMAP_14_53);
			MULT_54(13)<=signed(DIN_54_7)*signed(FMAP_14_54);
			MULT_55(13)<=signed(DIN_55_7)*signed(FMAP_14_55);
			MULT_56(13)<=signed(DIN_56_7)*signed(FMAP_14_56);
			MULT_57(13)<=signed(DIN_57_7)*signed(FMAP_14_57);
			MULT_58(13)<=signed(DIN_58_7)*signed(FMAP_14_58);
			MULT_59(13)<=signed(DIN_59_7)*signed(FMAP_14_59);
			MULT_60(13)<=signed(DIN_60_7)*signed(FMAP_14_60);
			MULT_61(13)<=signed(DIN_61_7)*signed(FMAP_14_61);
			MULT_62(13)<=signed(DIN_62_7)*signed(FMAP_14_62);
			MULT_63(13)<=signed(DIN_63_7)*signed(FMAP_14_63);
			MULT_64(13)<=signed(DIN_64_7)*signed(FMAP_14_64);
			MULT_65(13)<=signed(DIN_65_7)*signed(FMAP_14_65);
			MULT_66(13)<=signed(DIN_66_7)*signed(FMAP_14_66);
			MULT_67(13)<=signed(DIN_67_7)*signed(FMAP_14_67);
			MULT_68(13)<=signed(DIN_68_7)*signed(FMAP_14_68);
			MULT_69(13)<=signed(DIN_69_7)*signed(FMAP_14_69);
			MULT_70(13)<=signed(DIN_70_7)*signed(FMAP_14_70);
			MULT_71(13)<=signed(DIN_71_7)*signed(FMAP_14_71);
			MULT_72(13)<=signed(DIN_72_7)*signed(FMAP_14_72);
			MULT_73(13)<=signed(DIN_73_7)*signed(FMAP_14_73);
			MULT_74(13)<=signed(DIN_74_7)*signed(FMAP_14_74);
			MULT_75(13)<=signed(DIN_75_7)*signed(FMAP_14_75);
			MULT_76(13)<=signed(DIN_76_7)*signed(FMAP_14_76);
			MULT_77(13)<=signed(DIN_77_7)*signed(FMAP_14_77);
			MULT_78(13)<=signed(DIN_78_7)*signed(FMAP_14_78);
			MULT_79(13)<=signed(DIN_79_7)*signed(FMAP_14_79);
			MULT_80(13)<=signed(DIN_80_7)*signed(FMAP_14_80);
			MULT_81(13)<=signed(DIN_81_7)*signed(FMAP_14_81);
			MULT_82(13)<=signed(DIN_82_7)*signed(FMAP_14_82);
			MULT_83(13)<=signed(DIN_83_7)*signed(FMAP_14_83);
			MULT_84(13)<=signed(DIN_84_7)*signed(FMAP_14_84);
			MULT_85(13)<=signed(DIN_85_7)*signed(FMAP_14_85);
			MULT_86(13)<=signed(DIN_86_7)*signed(FMAP_14_86);
			MULT_87(13)<=signed(DIN_87_7)*signed(FMAP_14_87);
			MULT_88(13)<=signed(DIN_88_7)*signed(FMAP_14_88);
			MULT_89(13)<=signed(DIN_89_7)*signed(FMAP_14_89);
			MULT_90(13)<=signed(DIN_90_7)*signed(FMAP_14_90);
			MULT_91(13)<=signed(DIN_91_7)*signed(FMAP_14_91);
			MULT_92(13)<=signed(DIN_92_7)*signed(FMAP_14_92);
			MULT_93(13)<=signed(DIN_93_7)*signed(FMAP_14_93);
			MULT_94(13)<=signed(DIN_94_7)*signed(FMAP_14_94);
			MULT_95(13)<=signed(DIN_95_7)*signed(FMAP_14_95);
			MULT_96(13)<=signed(DIN_96_7)*signed(FMAP_14_96);
			MULT_97(13)<=signed(DIN_97_7)*signed(FMAP_14_97);
			MULT_98(13)<=signed(DIN_98_7)*signed(FMAP_14_98);
			MULT_99(13)<=signed(DIN_99_7)*signed(FMAP_14_99);
			MULT_100(13)<=signed(DIN_100_7)*signed(FMAP_14_100);
			MULT_101(13)<=signed(DIN_101_7)*signed(FMAP_14_101);
			MULT_102(13)<=signed(DIN_102_7)*signed(FMAP_14_102);
			MULT_103(13)<=signed(DIN_103_7)*signed(FMAP_14_103);
			MULT_104(13)<=signed(DIN_104_7)*signed(FMAP_14_104);
			MULT_105(13)<=signed(DIN_105_7)*signed(FMAP_14_105);
			MULT_106(13)<=signed(DIN_106_7)*signed(FMAP_14_106);
			MULT_107(13)<=signed(DIN_107_7)*signed(FMAP_14_107);
			MULT_108(13)<=signed(DIN_108_7)*signed(FMAP_14_108);
			MULT_109(13)<=signed(DIN_109_7)*signed(FMAP_14_109);
			MULT_110(13)<=signed(DIN_110_7)*signed(FMAP_14_110);
			MULT_111(13)<=signed(DIN_111_7)*signed(FMAP_14_111);
			MULT_112(13)<=signed(DIN_112_7)*signed(FMAP_14_112);
			MULT_113(13)<=signed(DIN_113_7)*signed(FMAP_14_113);
			MULT_114(13)<=signed(DIN_114_7)*signed(FMAP_14_114);
			MULT_115(13)<=signed(DIN_115_7)*signed(FMAP_14_115);
			MULT_116(13)<=signed(DIN_116_7)*signed(FMAP_14_116);
			MULT_117(13)<=signed(DIN_117_7)*signed(FMAP_14_117);
			MULT_118(13)<=signed(DIN_118_7)*signed(FMAP_14_118);
			MULT_119(13)<=signed(DIN_119_7)*signed(FMAP_14_119);
			MULT_120(13)<=signed(DIN_120_7)*signed(FMAP_14_120);

			MULT_1(14)<=signed(DIN_1_7)*signed(FMAP_15_1);
			MULT_2(14)<=signed(DIN_2_7)*signed(FMAP_15_2);
			MULT_3(14)<=signed(DIN_3_7)*signed(FMAP_15_3);
			MULT_4(14)<=signed(DIN_4_7)*signed(FMAP_15_4);
			MULT_5(14)<=signed(DIN_5_7)*signed(FMAP_15_5);
			MULT_6(14)<=signed(DIN_6_7)*signed(FMAP_15_6);
			MULT_7(14)<=signed(DIN_7_7)*signed(FMAP_15_7);
			MULT_8(14)<=signed(DIN_8_7)*signed(FMAP_15_8);
			MULT_9(14)<=signed(DIN_9_7)*signed(FMAP_15_9);
			MULT_10(14)<=signed(DIN_10_7)*signed(FMAP_15_10);
			MULT_11(14)<=signed(DIN_11_7)*signed(FMAP_15_11);
			MULT_12(14)<=signed(DIN_12_7)*signed(FMAP_15_12);
			MULT_13(14)<=signed(DIN_13_7)*signed(FMAP_15_13);
			MULT_14(14)<=signed(DIN_14_7)*signed(FMAP_15_14);
			MULT_15(14)<=signed(DIN_15_7)*signed(FMAP_15_15);
			MULT_16(14)<=signed(DIN_16_7)*signed(FMAP_15_16);
			MULT_17(14)<=signed(DIN_17_7)*signed(FMAP_15_17);
			MULT_18(14)<=signed(DIN_18_7)*signed(FMAP_15_18);
			MULT_19(14)<=signed(DIN_19_7)*signed(FMAP_15_19);
			MULT_20(14)<=signed(DIN_20_7)*signed(FMAP_15_20);
			MULT_21(14)<=signed(DIN_21_7)*signed(FMAP_15_21);
			MULT_22(14)<=signed(DIN_22_7)*signed(FMAP_15_22);
			MULT_23(14)<=signed(DIN_23_7)*signed(FMAP_15_23);
			MULT_24(14)<=signed(DIN_24_7)*signed(FMAP_15_24);
			MULT_25(14)<=signed(DIN_25_7)*signed(FMAP_15_25);
			MULT_26(14)<=signed(DIN_26_7)*signed(FMAP_15_26);
			MULT_27(14)<=signed(DIN_27_7)*signed(FMAP_15_27);
			MULT_28(14)<=signed(DIN_28_7)*signed(FMAP_15_28);
			MULT_29(14)<=signed(DIN_29_7)*signed(FMAP_15_29);
			MULT_30(14)<=signed(DIN_30_7)*signed(FMAP_15_30);
			MULT_31(14)<=signed(DIN_31_7)*signed(FMAP_15_31);
			MULT_32(14)<=signed(DIN_32_7)*signed(FMAP_15_32);
			MULT_33(14)<=signed(DIN_33_7)*signed(FMAP_15_33);
			MULT_34(14)<=signed(DIN_34_7)*signed(FMAP_15_34);
			MULT_35(14)<=signed(DIN_35_7)*signed(FMAP_15_35);
			MULT_36(14)<=signed(DIN_36_7)*signed(FMAP_15_36);
			MULT_37(14)<=signed(DIN_37_7)*signed(FMAP_15_37);
			MULT_38(14)<=signed(DIN_38_7)*signed(FMAP_15_38);
			MULT_39(14)<=signed(DIN_39_7)*signed(FMAP_15_39);
			MULT_40(14)<=signed(DIN_40_7)*signed(FMAP_15_40);
			MULT_41(14)<=signed(DIN_41_7)*signed(FMAP_15_41);
			MULT_42(14)<=signed(DIN_42_7)*signed(FMAP_15_42);
			MULT_43(14)<=signed(DIN_43_7)*signed(FMAP_15_43);
			MULT_44(14)<=signed(DIN_44_7)*signed(FMAP_15_44);
			MULT_45(14)<=signed(DIN_45_7)*signed(FMAP_15_45);
			MULT_46(14)<=signed(DIN_46_7)*signed(FMAP_15_46);
			MULT_47(14)<=signed(DIN_47_7)*signed(FMAP_15_47);
			MULT_48(14)<=signed(DIN_48_7)*signed(FMAP_15_48);
			MULT_49(14)<=signed(DIN_49_7)*signed(FMAP_15_49);
			MULT_50(14)<=signed(DIN_50_7)*signed(FMAP_15_50);
			MULT_51(14)<=signed(DIN_51_7)*signed(FMAP_15_51);
			MULT_52(14)<=signed(DIN_52_7)*signed(FMAP_15_52);
			MULT_53(14)<=signed(DIN_53_7)*signed(FMAP_15_53);
			MULT_54(14)<=signed(DIN_54_7)*signed(FMAP_15_54);
			MULT_55(14)<=signed(DIN_55_7)*signed(FMAP_15_55);
			MULT_56(14)<=signed(DIN_56_7)*signed(FMAP_15_56);
			MULT_57(14)<=signed(DIN_57_7)*signed(FMAP_15_57);
			MULT_58(14)<=signed(DIN_58_7)*signed(FMAP_15_58);
			MULT_59(14)<=signed(DIN_59_7)*signed(FMAP_15_59);
			MULT_60(14)<=signed(DIN_60_7)*signed(FMAP_15_60);
			MULT_61(14)<=signed(DIN_61_7)*signed(FMAP_15_61);
			MULT_62(14)<=signed(DIN_62_7)*signed(FMAP_15_62);
			MULT_63(14)<=signed(DIN_63_7)*signed(FMAP_15_63);
			MULT_64(14)<=signed(DIN_64_7)*signed(FMAP_15_64);
			MULT_65(14)<=signed(DIN_65_7)*signed(FMAP_15_65);
			MULT_66(14)<=signed(DIN_66_7)*signed(FMAP_15_66);
			MULT_67(14)<=signed(DIN_67_7)*signed(FMAP_15_67);
			MULT_68(14)<=signed(DIN_68_7)*signed(FMAP_15_68);
			MULT_69(14)<=signed(DIN_69_7)*signed(FMAP_15_69);
			MULT_70(14)<=signed(DIN_70_7)*signed(FMAP_15_70);
			MULT_71(14)<=signed(DIN_71_7)*signed(FMAP_15_71);
			MULT_72(14)<=signed(DIN_72_7)*signed(FMAP_15_72);
			MULT_73(14)<=signed(DIN_73_7)*signed(FMAP_15_73);
			MULT_74(14)<=signed(DIN_74_7)*signed(FMAP_15_74);
			MULT_75(14)<=signed(DIN_75_7)*signed(FMAP_15_75);
			MULT_76(14)<=signed(DIN_76_7)*signed(FMAP_15_76);
			MULT_77(14)<=signed(DIN_77_7)*signed(FMAP_15_77);
			MULT_78(14)<=signed(DIN_78_7)*signed(FMAP_15_78);
			MULT_79(14)<=signed(DIN_79_7)*signed(FMAP_15_79);
			MULT_80(14)<=signed(DIN_80_7)*signed(FMAP_15_80);
			MULT_81(14)<=signed(DIN_81_7)*signed(FMAP_15_81);
			MULT_82(14)<=signed(DIN_82_7)*signed(FMAP_15_82);
			MULT_83(14)<=signed(DIN_83_7)*signed(FMAP_15_83);
			MULT_84(14)<=signed(DIN_84_7)*signed(FMAP_15_84);
			MULT_85(14)<=signed(DIN_85_7)*signed(FMAP_15_85);
			MULT_86(14)<=signed(DIN_86_7)*signed(FMAP_15_86);
			MULT_87(14)<=signed(DIN_87_7)*signed(FMAP_15_87);
			MULT_88(14)<=signed(DIN_88_7)*signed(FMAP_15_88);
			MULT_89(14)<=signed(DIN_89_7)*signed(FMAP_15_89);
			MULT_90(14)<=signed(DIN_90_7)*signed(FMAP_15_90);
			MULT_91(14)<=signed(DIN_91_7)*signed(FMAP_15_91);
			MULT_92(14)<=signed(DIN_92_7)*signed(FMAP_15_92);
			MULT_93(14)<=signed(DIN_93_7)*signed(FMAP_15_93);
			MULT_94(14)<=signed(DIN_94_7)*signed(FMAP_15_94);
			MULT_95(14)<=signed(DIN_95_7)*signed(FMAP_15_95);
			MULT_96(14)<=signed(DIN_96_7)*signed(FMAP_15_96);
			MULT_97(14)<=signed(DIN_97_7)*signed(FMAP_15_97);
			MULT_98(14)<=signed(DIN_98_7)*signed(FMAP_15_98);
			MULT_99(14)<=signed(DIN_99_7)*signed(FMAP_15_99);
			MULT_100(14)<=signed(DIN_100_7)*signed(FMAP_15_100);
			MULT_101(14)<=signed(DIN_101_7)*signed(FMAP_15_101);
			MULT_102(14)<=signed(DIN_102_7)*signed(FMAP_15_102);
			MULT_103(14)<=signed(DIN_103_7)*signed(FMAP_15_103);
			MULT_104(14)<=signed(DIN_104_7)*signed(FMAP_15_104);
			MULT_105(14)<=signed(DIN_105_7)*signed(FMAP_15_105);
			MULT_106(14)<=signed(DIN_106_7)*signed(FMAP_15_106);
			MULT_107(14)<=signed(DIN_107_7)*signed(FMAP_15_107);
			MULT_108(14)<=signed(DIN_108_7)*signed(FMAP_15_108);
			MULT_109(14)<=signed(DIN_109_7)*signed(FMAP_15_109);
			MULT_110(14)<=signed(DIN_110_7)*signed(FMAP_15_110);
			MULT_111(14)<=signed(DIN_111_7)*signed(FMAP_15_111);
			MULT_112(14)<=signed(DIN_112_7)*signed(FMAP_15_112);
			MULT_113(14)<=signed(DIN_113_7)*signed(FMAP_15_113);
			MULT_114(14)<=signed(DIN_114_7)*signed(FMAP_15_114);
			MULT_115(14)<=signed(DIN_115_7)*signed(FMAP_15_115);
			MULT_116(14)<=signed(DIN_116_7)*signed(FMAP_15_116);
			MULT_117(14)<=signed(DIN_117_7)*signed(FMAP_15_117);
			MULT_118(14)<=signed(DIN_118_7)*signed(FMAP_15_118);
			MULT_119(14)<=signed(DIN_119_7)*signed(FMAP_15_119);
			MULT_120(14)<=signed(DIN_120_7)*signed(FMAP_15_120);

			MULT_1(15)<=signed(DIN_1_7)*signed(FMAP_16_1);
			MULT_2(15)<=signed(DIN_2_7)*signed(FMAP_16_2);
			MULT_3(15)<=signed(DIN_3_7)*signed(FMAP_16_3);
			MULT_4(15)<=signed(DIN_4_7)*signed(FMAP_16_4);
			MULT_5(15)<=signed(DIN_5_7)*signed(FMAP_16_5);
			MULT_6(15)<=signed(DIN_6_7)*signed(FMAP_16_6);
			MULT_7(15)<=signed(DIN_7_7)*signed(FMAP_16_7);
			MULT_8(15)<=signed(DIN_8_7)*signed(FMAP_16_8);
			MULT_9(15)<=signed(DIN_9_7)*signed(FMAP_16_9);
			MULT_10(15)<=signed(DIN_10_7)*signed(FMAP_16_10);
			MULT_11(15)<=signed(DIN_11_7)*signed(FMAP_16_11);
			MULT_12(15)<=signed(DIN_12_7)*signed(FMAP_16_12);
			MULT_13(15)<=signed(DIN_13_7)*signed(FMAP_16_13);
			MULT_14(15)<=signed(DIN_14_7)*signed(FMAP_16_14);
			MULT_15(15)<=signed(DIN_15_7)*signed(FMAP_16_15);
			MULT_16(15)<=signed(DIN_16_7)*signed(FMAP_16_16);
			MULT_17(15)<=signed(DIN_17_7)*signed(FMAP_16_17);
			MULT_18(15)<=signed(DIN_18_7)*signed(FMAP_16_18);
			MULT_19(15)<=signed(DIN_19_7)*signed(FMAP_16_19);
			MULT_20(15)<=signed(DIN_20_7)*signed(FMAP_16_20);
			MULT_21(15)<=signed(DIN_21_7)*signed(FMAP_16_21);
			MULT_22(15)<=signed(DIN_22_7)*signed(FMAP_16_22);
			MULT_23(15)<=signed(DIN_23_7)*signed(FMAP_16_23);
			MULT_24(15)<=signed(DIN_24_7)*signed(FMAP_16_24);
			MULT_25(15)<=signed(DIN_25_7)*signed(FMAP_16_25);
			MULT_26(15)<=signed(DIN_26_7)*signed(FMAP_16_26);
			MULT_27(15)<=signed(DIN_27_7)*signed(FMAP_16_27);
			MULT_28(15)<=signed(DIN_28_7)*signed(FMAP_16_28);
			MULT_29(15)<=signed(DIN_29_7)*signed(FMAP_16_29);
			MULT_30(15)<=signed(DIN_30_7)*signed(FMAP_16_30);
			MULT_31(15)<=signed(DIN_31_7)*signed(FMAP_16_31);
			MULT_32(15)<=signed(DIN_32_7)*signed(FMAP_16_32);
			MULT_33(15)<=signed(DIN_33_7)*signed(FMAP_16_33);
			MULT_34(15)<=signed(DIN_34_7)*signed(FMAP_16_34);
			MULT_35(15)<=signed(DIN_35_7)*signed(FMAP_16_35);
			MULT_36(15)<=signed(DIN_36_7)*signed(FMAP_16_36);
			MULT_37(15)<=signed(DIN_37_7)*signed(FMAP_16_37);
			MULT_38(15)<=signed(DIN_38_7)*signed(FMAP_16_38);
			MULT_39(15)<=signed(DIN_39_7)*signed(FMAP_16_39);
			MULT_40(15)<=signed(DIN_40_7)*signed(FMAP_16_40);
			MULT_41(15)<=signed(DIN_41_7)*signed(FMAP_16_41);
			MULT_42(15)<=signed(DIN_42_7)*signed(FMAP_16_42);
			MULT_43(15)<=signed(DIN_43_7)*signed(FMAP_16_43);
			MULT_44(15)<=signed(DIN_44_7)*signed(FMAP_16_44);
			MULT_45(15)<=signed(DIN_45_7)*signed(FMAP_16_45);
			MULT_46(15)<=signed(DIN_46_7)*signed(FMAP_16_46);
			MULT_47(15)<=signed(DIN_47_7)*signed(FMAP_16_47);
			MULT_48(15)<=signed(DIN_48_7)*signed(FMAP_16_48);
			MULT_49(15)<=signed(DIN_49_7)*signed(FMAP_16_49);
			MULT_50(15)<=signed(DIN_50_7)*signed(FMAP_16_50);
			MULT_51(15)<=signed(DIN_51_7)*signed(FMAP_16_51);
			MULT_52(15)<=signed(DIN_52_7)*signed(FMAP_16_52);
			MULT_53(15)<=signed(DIN_53_7)*signed(FMAP_16_53);
			MULT_54(15)<=signed(DIN_54_7)*signed(FMAP_16_54);
			MULT_55(15)<=signed(DIN_55_7)*signed(FMAP_16_55);
			MULT_56(15)<=signed(DIN_56_7)*signed(FMAP_16_56);
			MULT_57(15)<=signed(DIN_57_7)*signed(FMAP_16_57);
			MULT_58(15)<=signed(DIN_58_7)*signed(FMAP_16_58);
			MULT_59(15)<=signed(DIN_59_7)*signed(FMAP_16_59);
			MULT_60(15)<=signed(DIN_60_7)*signed(FMAP_16_60);
			MULT_61(15)<=signed(DIN_61_7)*signed(FMAP_16_61);
			MULT_62(15)<=signed(DIN_62_7)*signed(FMAP_16_62);
			MULT_63(15)<=signed(DIN_63_7)*signed(FMAP_16_63);
			MULT_64(15)<=signed(DIN_64_7)*signed(FMAP_16_64);
			MULT_65(15)<=signed(DIN_65_7)*signed(FMAP_16_65);
			MULT_66(15)<=signed(DIN_66_7)*signed(FMAP_16_66);
			MULT_67(15)<=signed(DIN_67_7)*signed(FMAP_16_67);
			MULT_68(15)<=signed(DIN_68_7)*signed(FMAP_16_68);
			MULT_69(15)<=signed(DIN_69_7)*signed(FMAP_16_69);
			MULT_70(15)<=signed(DIN_70_7)*signed(FMAP_16_70);
			MULT_71(15)<=signed(DIN_71_7)*signed(FMAP_16_71);
			MULT_72(15)<=signed(DIN_72_7)*signed(FMAP_16_72);
			MULT_73(15)<=signed(DIN_73_7)*signed(FMAP_16_73);
			MULT_74(15)<=signed(DIN_74_7)*signed(FMAP_16_74);
			MULT_75(15)<=signed(DIN_75_7)*signed(FMAP_16_75);
			MULT_76(15)<=signed(DIN_76_7)*signed(FMAP_16_76);
			MULT_77(15)<=signed(DIN_77_7)*signed(FMAP_16_77);
			MULT_78(15)<=signed(DIN_78_7)*signed(FMAP_16_78);
			MULT_79(15)<=signed(DIN_79_7)*signed(FMAP_16_79);
			MULT_80(15)<=signed(DIN_80_7)*signed(FMAP_16_80);
			MULT_81(15)<=signed(DIN_81_7)*signed(FMAP_16_81);
			MULT_82(15)<=signed(DIN_82_7)*signed(FMAP_16_82);
			MULT_83(15)<=signed(DIN_83_7)*signed(FMAP_16_83);
			MULT_84(15)<=signed(DIN_84_7)*signed(FMAP_16_84);
			MULT_85(15)<=signed(DIN_85_7)*signed(FMAP_16_85);
			MULT_86(15)<=signed(DIN_86_7)*signed(FMAP_16_86);
			MULT_87(15)<=signed(DIN_87_7)*signed(FMAP_16_87);
			MULT_88(15)<=signed(DIN_88_7)*signed(FMAP_16_88);
			MULT_89(15)<=signed(DIN_89_7)*signed(FMAP_16_89);
			MULT_90(15)<=signed(DIN_90_7)*signed(FMAP_16_90);
			MULT_91(15)<=signed(DIN_91_7)*signed(FMAP_16_91);
			MULT_92(15)<=signed(DIN_92_7)*signed(FMAP_16_92);
			MULT_93(15)<=signed(DIN_93_7)*signed(FMAP_16_93);
			MULT_94(15)<=signed(DIN_94_7)*signed(FMAP_16_94);
			MULT_95(15)<=signed(DIN_95_7)*signed(FMAP_16_95);
			MULT_96(15)<=signed(DIN_96_7)*signed(FMAP_16_96);
			MULT_97(15)<=signed(DIN_97_7)*signed(FMAP_16_97);
			MULT_98(15)<=signed(DIN_98_7)*signed(FMAP_16_98);
			MULT_99(15)<=signed(DIN_99_7)*signed(FMAP_16_99);
			MULT_100(15)<=signed(DIN_100_7)*signed(FMAP_16_100);
			MULT_101(15)<=signed(DIN_101_7)*signed(FMAP_16_101);
			MULT_102(15)<=signed(DIN_102_7)*signed(FMAP_16_102);
			MULT_103(15)<=signed(DIN_103_7)*signed(FMAP_16_103);
			MULT_104(15)<=signed(DIN_104_7)*signed(FMAP_16_104);
			MULT_105(15)<=signed(DIN_105_7)*signed(FMAP_16_105);
			MULT_106(15)<=signed(DIN_106_7)*signed(FMAP_16_106);
			MULT_107(15)<=signed(DIN_107_7)*signed(FMAP_16_107);
			MULT_108(15)<=signed(DIN_108_7)*signed(FMAP_16_108);
			MULT_109(15)<=signed(DIN_109_7)*signed(FMAP_16_109);
			MULT_110(15)<=signed(DIN_110_7)*signed(FMAP_16_110);
			MULT_111(15)<=signed(DIN_111_7)*signed(FMAP_16_111);
			MULT_112(15)<=signed(DIN_112_7)*signed(FMAP_16_112);
			MULT_113(15)<=signed(DIN_113_7)*signed(FMAP_16_113);
			MULT_114(15)<=signed(DIN_114_7)*signed(FMAP_16_114);
			MULT_115(15)<=signed(DIN_115_7)*signed(FMAP_16_115);
			MULT_116(15)<=signed(DIN_116_7)*signed(FMAP_16_116);
			MULT_117(15)<=signed(DIN_117_7)*signed(FMAP_16_117);
			MULT_118(15)<=signed(DIN_118_7)*signed(FMAP_16_118);
			MULT_119(15)<=signed(DIN_119_7)*signed(FMAP_16_119);
			MULT_120(15)<=signed(DIN_120_7)*signed(FMAP_16_120);

			MULT_1(16)<=signed(DIN_1_7)*signed(FMAP_17_1);
			MULT_2(16)<=signed(DIN_2_7)*signed(FMAP_17_2);
			MULT_3(16)<=signed(DIN_3_7)*signed(FMAP_17_3);
			MULT_4(16)<=signed(DIN_4_7)*signed(FMAP_17_4);
			MULT_5(16)<=signed(DIN_5_7)*signed(FMAP_17_5);
			MULT_6(16)<=signed(DIN_6_7)*signed(FMAP_17_6);
			MULT_7(16)<=signed(DIN_7_7)*signed(FMAP_17_7);
			MULT_8(16)<=signed(DIN_8_7)*signed(FMAP_17_8);
			MULT_9(16)<=signed(DIN_9_7)*signed(FMAP_17_9);
			MULT_10(16)<=signed(DIN_10_7)*signed(FMAP_17_10);
			MULT_11(16)<=signed(DIN_11_7)*signed(FMAP_17_11);
			MULT_12(16)<=signed(DIN_12_7)*signed(FMAP_17_12);
			MULT_13(16)<=signed(DIN_13_7)*signed(FMAP_17_13);
			MULT_14(16)<=signed(DIN_14_7)*signed(FMAP_17_14);
			MULT_15(16)<=signed(DIN_15_7)*signed(FMAP_17_15);
			MULT_16(16)<=signed(DIN_16_7)*signed(FMAP_17_16);
			MULT_17(16)<=signed(DIN_17_7)*signed(FMAP_17_17);
			MULT_18(16)<=signed(DIN_18_7)*signed(FMAP_17_18);
			MULT_19(16)<=signed(DIN_19_7)*signed(FMAP_17_19);
			MULT_20(16)<=signed(DIN_20_7)*signed(FMAP_17_20);
			MULT_21(16)<=signed(DIN_21_7)*signed(FMAP_17_21);
			MULT_22(16)<=signed(DIN_22_7)*signed(FMAP_17_22);
			MULT_23(16)<=signed(DIN_23_7)*signed(FMAP_17_23);
			MULT_24(16)<=signed(DIN_24_7)*signed(FMAP_17_24);
			MULT_25(16)<=signed(DIN_25_7)*signed(FMAP_17_25);
			MULT_26(16)<=signed(DIN_26_7)*signed(FMAP_17_26);
			MULT_27(16)<=signed(DIN_27_7)*signed(FMAP_17_27);
			MULT_28(16)<=signed(DIN_28_7)*signed(FMAP_17_28);
			MULT_29(16)<=signed(DIN_29_7)*signed(FMAP_17_29);
			MULT_30(16)<=signed(DIN_30_7)*signed(FMAP_17_30);
			MULT_31(16)<=signed(DIN_31_7)*signed(FMAP_17_31);
			MULT_32(16)<=signed(DIN_32_7)*signed(FMAP_17_32);
			MULT_33(16)<=signed(DIN_33_7)*signed(FMAP_17_33);
			MULT_34(16)<=signed(DIN_34_7)*signed(FMAP_17_34);
			MULT_35(16)<=signed(DIN_35_7)*signed(FMAP_17_35);
			MULT_36(16)<=signed(DIN_36_7)*signed(FMAP_17_36);
			MULT_37(16)<=signed(DIN_37_7)*signed(FMAP_17_37);
			MULT_38(16)<=signed(DIN_38_7)*signed(FMAP_17_38);
			MULT_39(16)<=signed(DIN_39_7)*signed(FMAP_17_39);
			MULT_40(16)<=signed(DIN_40_7)*signed(FMAP_17_40);
			MULT_41(16)<=signed(DIN_41_7)*signed(FMAP_17_41);
			MULT_42(16)<=signed(DIN_42_7)*signed(FMAP_17_42);
			MULT_43(16)<=signed(DIN_43_7)*signed(FMAP_17_43);
			MULT_44(16)<=signed(DIN_44_7)*signed(FMAP_17_44);
			MULT_45(16)<=signed(DIN_45_7)*signed(FMAP_17_45);
			MULT_46(16)<=signed(DIN_46_7)*signed(FMAP_17_46);
			MULT_47(16)<=signed(DIN_47_7)*signed(FMAP_17_47);
			MULT_48(16)<=signed(DIN_48_7)*signed(FMAP_17_48);
			MULT_49(16)<=signed(DIN_49_7)*signed(FMAP_17_49);
			MULT_50(16)<=signed(DIN_50_7)*signed(FMAP_17_50);
			MULT_51(16)<=signed(DIN_51_7)*signed(FMAP_17_51);
			MULT_52(16)<=signed(DIN_52_7)*signed(FMAP_17_52);
			MULT_53(16)<=signed(DIN_53_7)*signed(FMAP_17_53);
			MULT_54(16)<=signed(DIN_54_7)*signed(FMAP_17_54);
			MULT_55(16)<=signed(DIN_55_7)*signed(FMAP_17_55);
			MULT_56(16)<=signed(DIN_56_7)*signed(FMAP_17_56);
			MULT_57(16)<=signed(DIN_57_7)*signed(FMAP_17_57);
			MULT_58(16)<=signed(DIN_58_7)*signed(FMAP_17_58);
			MULT_59(16)<=signed(DIN_59_7)*signed(FMAP_17_59);
			MULT_60(16)<=signed(DIN_60_7)*signed(FMAP_17_60);
			MULT_61(16)<=signed(DIN_61_7)*signed(FMAP_17_61);
			MULT_62(16)<=signed(DIN_62_7)*signed(FMAP_17_62);
			MULT_63(16)<=signed(DIN_63_7)*signed(FMAP_17_63);
			MULT_64(16)<=signed(DIN_64_7)*signed(FMAP_17_64);
			MULT_65(16)<=signed(DIN_65_7)*signed(FMAP_17_65);
			MULT_66(16)<=signed(DIN_66_7)*signed(FMAP_17_66);
			MULT_67(16)<=signed(DIN_67_7)*signed(FMAP_17_67);
			MULT_68(16)<=signed(DIN_68_7)*signed(FMAP_17_68);
			MULT_69(16)<=signed(DIN_69_7)*signed(FMAP_17_69);
			MULT_70(16)<=signed(DIN_70_7)*signed(FMAP_17_70);
			MULT_71(16)<=signed(DIN_71_7)*signed(FMAP_17_71);
			MULT_72(16)<=signed(DIN_72_7)*signed(FMAP_17_72);
			MULT_73(16)<=signed(DIN_73_7)*signed(FMAP_17_73);
			MULT_74(16)<=signed(DIN_74_7)*signed(FMAP_17_74);
			MULT_75(16)<=signed(DIN_75_7)*signed(FMAP_17_75);
			MULT_76(16)<=signed(DIN_76_7)*signed(FMAP_17_76);
			MULT_77(16)<=signed(DIN_77_7)*signed(FMAP_17_77);
			MULT_78(16)<=signed(DIN_78_7)*signed(FMAP_17_78);
			MULT_79(16)<=signed(DIN_79_7)*signed(FMAP_17_79);
			MULT_80(16)<=signed(DIN_80_7)*signed(FMAP_17_80);
			MULT_81(16)<=signed(DIN_81_7)*signed(FMAP_17_81);
			MULT_82(16)<=signed(DIN_82_7)*signed(FMAP_17_82);
			MULT_83(16)<=signed(DIN_83_7)*signed(FMAP_17_83);
			MULT_84(16)<=signed(DIN_84_7)*signed(FMAP_17_84);
			MULT_85(16)<=signed(DIN_85_7)*signed(FMAP_17_85);
			MULT_86(16)<=signed(DIN_86_7)*signed(FMAP_17_86);
			MULT_87(16)<=signed(DIN_87_7)*signed(FMAP_17_87);
			MULT_88(16)<=signed(DIN_88_7)*signed(FMAP_17_88);
			MULT_89(16)<=signed(DIN_89_7)*signed(FMAP_17_89);
			MULT_90(16)<=signed(DIN_90_7)*signed(FMAP_17_90);
			MULT_91(16)<=signed(DIN_91_7)*signed(FMAP_17_91);
			MULT_92(16)<=signed(DIN_92_7)*signed(FMAP_17_92);
			MULT_93(16)<=signed(DIN_93_7)*signed(FMAP_17_93);
			MULT_94(16)<=signed(DIN_94_7)*signed(FMAP_17_94);
			MULT_95(16)<=signed(DIN_95_7)*signed(FMAP_17_95);
			MULT_96(16)<=signed(DIN_96_7)*signed(FMAP_17_96);
			MULT_97(16)<=signed(DIN_97_7)*signed(FMAP_17_97);
			MULT_98(16)<=signed(DIN_98_7)*signed(FMAP_17_98);
			MULT_99(16)<=signed(DIN_99_7)*signed(FMAP_17_99);
			MULT_100(16)<=signed(DIN_100_7)*signed(FMAP_17_100);
			MULT_101(16)<=signed(DIN_101_7)*signed(FMAP_17_101);
			MULT_102(16)<=signed(DIN_102_7)*signed(FMAP_17_102);
			MULT_103(16)<=signed(DIN_103_7)*signed(FMAP_17_103);
			MULT_104(16)<=signed(DIN_104_7)*signed(FMAP_17_104);
			MULT_105(16)<=signed(DIN_105_7)*signed(FMAP_17_105);
			MULT_106(16)<=signed(DIN_106_7)*signed(FMAP_17_106);
			MULT_107(16)<=signed(DIN_107_7)*signed(FMAP_17_107);
			MULT_108(16)<=signed(DIN_108_7)*signed(FMAP_17_108);
			MULT_109(16)<=signed(DIN_109_7)*signed(FMAP_17_109);
			MULT_110(16)<=signed(DIN_110_7)*signed(FMAP_17_110);
			MULT_111(16)<=signed(DIN_111_7)*signed(FMAP_17_111);
			MULT_112(16)<=signed(DIN_112_7)*signed(FMAP_17_112);
			MULT_113(16)<=signed(DIN_113_7)*signed(FMAP_17_113);
			MULT_114(16)<=signed(DIN_114_7)*signed(FMAP_17_114);
			MULT_115(16)<=signed(DIN_115_7)*signed(FMAP_17_115);
			MULT_116(16)<=signed(DIN_116_7)*signed(FMAP_17_116);
			MULT_117(16)<=signed(DIN_117_7)*signed(FMAP_17_117);
			MULT_118(16)<=signed(DIN_118_7)*signed(FMAP_17_118);
			MULT_119(16)<=signed(DIN_119_7)*signed(FMAP_17_119);
			MULT_120(16)<=signed(DIN_120_7)*signed(FMAP_17_120);

			MULT_1(17)<=signed(DIN_1_7)*signed(FMAP_18_1);
			MULT_2(17)<=signed(DIN_2_7)*signed(FMAP_18_2);
			MULT_3(17)<=signed(DIN_3_7)*signed(FMAP_18_3);
			MULT_4(17)<=signed(DIN_4_7)*signed(FMAP_18_4);
			MULT_5(17)<=signed(DIN_5_7)*signed(FMAP_18_5);
			MULT_6(17)<=signed(DIN_6_7)*signed(FMAP_18_6);
			MULT_7(17)<=signed(DIN_7_7)*signed(FMAP_18_7);
			MULT_8(17)<=signed(DIN_8_7)*signed(FMAP_18_8);
			MULT_9(17)<=signed(DIN_9_7)*signed(FMAP_18_9);
			MULT_10(17)<=signed(DIN_10_7)*signed(FMAP_18_10);
			MULT_11(17)<=signed(DIN_11_7)*signed(FMAP_18_11);
			MULT_12(17)<=signed(DIN_12_7)*signed(FMAP_18_12);
			MULT_13(17)<=signed(DIN_13_7)*signed(FMAP_18_13);
			MULT_14(17)<=signed(DIN_14_7)*signed(FMAP_18_14);
			MULT_15(17)<=signed(DIN_15_7)*signed(FMAP_18_15);
			MULT_16(17)<=signed(DIN_16_7)*signed(FMAP_18_16);
			MULT_17(17)<=signed(DIN_17_7)*signed(FMAP_18_17);
			MULT_18(17)<=signed(DIN_18_7)*signed(FMAP_18_18);
			MULT_19(17)<=signed(DIN_19_7)*signed(FMAP_18_19);
			MULT_20(17)<=signed(DIN_20_7)*signed(FMAP_18_20);
			MULT_21(17)<=signed(DIN_21_7)*signed(FMAP_18_21);
			MULT_22(17)<=signed(DIN_22_7)*signed(FMAP_18_22);
			MULT_23(17)<=signed(DIN_23_7)*signed(FMAP_18_23);
			MULT_24(17)<=signed(DIN_24_7)*signed(FMAP_18_24);
			MULT_25(17)<=signed(DIN_25_7)*signed(FMAP_18_25);
			MULT_26(17)<=signed(DIN_26_7)*signed(FMAP_18_26);
			MULT_27(17)<=signed(DIN_27_7)*signed(FMAP_18_27);
			MULT_28(17)<=signed(DIN_28_7)*signed(FMAP_18_28);
			MULT_29(17)<=signed(DIN_29_7)*signed(FMAP_18_29);
			MULT_30(17)<=signed(DIN_30_7)*signed(FMAP_18_30);
			MULT_31(17)<=signed(DIN_31_7)*signed(FMAP_18_31);
			MULT_32(17)<=signed(DIN_32_7)*signed(FMAP_18_32);
			MULT_33(17)<=signed(DIN_33_7)*signed(FMAP_18_33);
			MULT_34(17)<=signed(DIN_34_7)*signed(FMAP_18_34);
			MULT_35(17)<=signed(DIN_35_7)*signed(FMAP_18_35);
			MULT_36(17)<=signed(DIN_36_7)*signed(FMAP_18_36);
			MULT_37(17)<=signed(DIN_37_7)*signed(FMAP_18_37);
			MULT_38(17)<=signed(DIN_38_7)*signed(FMAP_18_38);
			MULT_39(17)<=signed(DIN_39_7)*signed(FMAP_18_39);
			MULT_40(17)<=signed(DIN_40_7)*signed(FMAP_18_40);
			MULT_41(17)<=signed(DIN_41_7)*signed(FMAP_18_41);
			MULT_42(17)<=signed(DIN_42_7)*signed(FMAP_18_42);
			MULT_43(17)<=signed(DIN_43_7)*signed(FMAP_18_43);
			MULT_44(17)<=signed(DIN_44_7)*signed(FMAP_18_44);
			MULT_45(17)<=signed(DIN_45_7)*signed(FMAP_18_45);
			MULT_46(17)<=signed(DIN_46_7)*signed(FMAP_18_46);
			MULT_47(17)<=signed(DIN_47_7)*signed(FMAP_18_47);
			MULT_48(17)<=signed(DIN_48_7)*signed(FMAP_18_48);
			MULT_49(17)<=signed(DIN_49_7)*signed(FMAP_18_49);
			MULT_50(17)<=signed(DIN_50_7)*signed(FMAP_18_50);
			MULT_51(17)<=signed(DIN_51_7)*signed(FMAP_18_51);
			MULT_52(17)<=signed(DIN_52_7)*signed(FMAP_18_52);
			MULT_53(17)<=signed(DIN_53_7)*signed(FMAP_18_53);
			MULT_54(17)<=signed(DIN_54_7)*signed(FMAP_18_54);
			MULT_55(17)<=signed(DIN_55_7)*signed(FMAP_18_55);
			MULT_56(17)<=signed(DIN_56_7)*signed(FMAP_18_56);
			MULT_57(17)<=signed(DIN_57_7)*signed(FMAP_18_57);
			MULT_58(17)<=signed(DIN_58_7)*signed(FMAP_18_58);
			MULT_59(17)<=signed(DIN_59_7)*signed(FMAP_18_59);
			MULT_60(17)<=signed(DIN_60_7)*signed(FMAP_18_60);
			MULT_61(17)<=signed(DIN_61_7)*signed(FMAP_18_61);
			MULT_62(17)<=signed(DIN_62_7)*signed(FMAP_18_62);
			MULT_63(17)<=signed(DIN_63_7)*signed(FMAP_18_63);
			MULT_64(17)<=signed(DIN_64_7)*signed(FMAP_18_64);
			MULT_65(17)<=signed(DIN_65_7)*signed(FMAP_18_65);
			MULT_66(17)<=signed(DIN_66_7)*signed(FMAP_18_66);
			MULT_67(17)<=signed(DIN_67_7)*signed(FMAP_18_67);
			MULT_68(17)<=signed(DIN_68_7)*signed(FMAP_18_68);
			MULT_69(17)<=signed(DIN_69_7)*signed(FMAP_18_69);
			MULT_70(17)<=signed(DIN_70_7)*signed(FMAP_18_70);
			MULT_71(17)<=signed(DIN_71_7)*signed(FMAP_18_71);
			MULT_72(17)<=signed(DIN_72_7)*signed(FMAP_18_72);
			MULT_73(17)<=signed(DIN_73_7)*signed(FMAP_18_73);
			MULT_74(17)<=signed(DIN_74_7)*signed(FMAP_18_74);
			MULT_75(17)<=signed(DIN_75_7)*signed(FMAP_18_75);
			MULT_76(17)<=signed(DIN_76_7)*signed(FMAP_18_76);
			MULT_77(17)<=signed(DIN_77_7)*signed(FMAP_18_77);
			MULT_78(17)<=signed(DIN_78_7)*signed(FMAP_18_78);
			MULT_79(17)<=signed(DIN_79_7)*signed(FMAP_18_79);
			MULT_80(17)<=signed(DIN_80_7)*signed(FMAP_18_80);
			MULT_81(17)<=signed(DIN_81_7)*signed(FMAP_18_81);
			MULT_82(17)<=signed(DIN_82_7)*signed(FMAP_18_82);
			MULT_83(17)<=signed(DIN_83_7)*signed(FMAP_18_83);
			MULT_84(17)<=signed(DIN_84_7)*signed(FMAP_18_84);
			MULT_85(17)<=signed(DIN_85_7)*signed(FMAP_18_85);
			MULT_86(17)<=signed(DIN_86_7)*signed(FMAP_18_86);
			MULT_87(17)<=signed(DIN_87_7)*signed(FMAP_18_87);
			MULT_88(17)<=signed(DIN_88_7)*signed(FMAP_18_88);
			MULT_89(17)<=signed(DIN_89_7)*signed(FMAP_18_89);
			MULT_90(17)<=signed(DIN_90_7)*signed(FMAP_18_90);
			MULT_91(17)<=signed(DIN_91_7)*signed(FMAP_18_91);
			MULT_92(17)<=signed(DIN_92_7)*signed(FMAP_18_92);
			MULT_93(17)<=signed(DIN_93_7)*signed(FMAP_18_93);
			MULT_94(17)<=signed(DIN_94_7)*signed(FMAP_18_94);
			MULT_95(17)<=signed(DIN_95_7)*signed(FMAP_18_95);
			MULT_96(17)<=signed(DIN_96_7)*signed(FMAP_18_96);
			MULT_97(17)<=signed(DIN_97_7)*signed(FMAP_18_97);
			MULT_98(17)<=signed(DIN_98_7)*signed(FMAP_18_98);
			MULT_99(17)<=signed(DIN_99_7)*signed(FMAP_18_99);
			MULT_100(17)<=signed(DIN_100_7)*signed(FMAP_18_100);
			MULT_101(17)<=signed(DIN_101_7)*signed(FMAP_18_101);
			MULT_102(17)<=signed(DIN_102_7)*signed(FMAP_18_102);
			MULT_103(17)<=signed(DIN_103_7)*signed(FMAP_18_103);
			MULT_104(17)<=signed(DIN_104_7)*signed(FMAP_18_104);
			MULT_105(17)<=signed(DIN_105_7)*signed(FMAP_18_105);
			MULT_106(17)<=signed(DIN_106_7)*signed(FMAP_18_106);
			MULT_107(17)<=signed(DIN_107_7)*signed(FMAP_18_107);
			MULT_108(17)<=signed(DIN_108_7)*signed(FMAP_18_108);
			MULT_109(17)<=signed(DIN_109_7)*signed(FMAP_18_109);
			MULT_110(17)<=signed(DIN_110_7)*signed(FMAP_18_110);
			MULT_111(17)<=signed(DIN_111_7)*signed(FMAP_18_111);
			MULT_112(17)<=signed(DIN_112_7)*signed(FMAP_18_112);
			MULT_113(17)<=signed(DIN_113_7)*signed(FMAP_18_113);
			MULT_114(17)<=signed(DIN_114_7)*signed(FMAP_18_114);
			MULT_115(17)<=signed(DIN_115_7)*signed(FMAP_18_115);
			MULT_116(17)<=signed(DIN_116_7)*signed(FMAP_18_116);
			MULT_117(17)<=signed(DIN_117_7)*signed(FMAP_18_117);
			MULT_118(17)<=signed(DIN_118_7)*signed(FMAP_18_118);
			MULT_119(17)<=signed(DIN_119_7)*signed(FMAP_18_119);
			MULT_120(17)<=signed(DIN_120_7)*signed(FMAP_18_120);

			MULT_1(18)<=signed(DIN_1_7)*signed(FMAP_19_1);
			MULT_2(18)<=signed(DIN_2_7)*signed(FMAP_19_2);
			MULT_3(18)<=signed(DIN_3_7)*signed(FMAP_19_3);
			MULT_4(18)<=signed(DIN_4_7)*signed(FMAP_19_4);
			MULT_5(18)<=signed(DIN_5_7)*signed(FMAP_19_5);
			MULT_6(18)<=signed(DIN_6_7)*signed(FMAP_19_6);
			MULT_7(18)<=signed(DIN_7_7)*signed(FMAP_19_7);
			MULT_8(18)<=signed(DIN_8_7)*signed(FMAP_19_8);
			MULT_9(18)<=signed(DIN_9_7)*signed(FMAP_19_9);
			MULT_10(18)<=signed(DIN_10_7)*signed(FMAP_19_10);
			MULT_11(18)<=signed(DIN_11_7)*signed(FMAP_19_11);
			MULT_12(18)<=signed(DIN_12_7)*signed(FMAP_19_12);
			MULT_13(18)<=signed(DIN_13_7)*signed(FMAP_19_13);
			MULT_14(18)<=signed(DIN_14_7)*signed(FMAP_19_14);
			MULT_15(18)<=signed(DIN_15_7)*signed(FMAP_19_15);
			MULT_16(18)<=signed(DIN_16_7)*signed(FMAP_19_16);
			MULT_17(18)<=signed(DIN_17_7)*signed(FMAP_19_17);
			MULT_18(18)<=signed(DIN_18_7)*signed(FMAP_19_18);
			MULT_19(18)<=signed(DIN_19_7)*signed(FMAP_19_19);
			MULT_20(18)<=signed(DIN_20_7)*signed(FMAP_19_20);
			MULT_21(18)<=signed(DIN_21_7)*signed(FMAP_19_21);
			MULT_22(18)<=signed(DIN_22_7)*signed(FMAP_19_22);
			MULT_23(18)<=signed(DIN_23_7)*signed(FMAP_19_23);
			MULT_24(18)<=signed(DIN_24_7)*signed(FMAP_19_24);
			MULT_25(18)<=signed(DIN_25_7)*signed(FMAP_19_25);
			MULT_26(18)<=signed(DIN_26_7)*signed(FMAP_19_26);
			MULT_27(18)<=signed(DIN_27_7)*signed(FMAP_19_27);
			MULT_28(18)<=signed(DIN_28_7)*signed(FMAP_19_28);
			MULT_29(18)<=signed(DIN_29_7)*signed(FMAP_19_29);
			MULT_30(18)<=signed(DIN_30_7)*signed(FMAP_19_30);
			MULT_31(18)<=signed(DIN_31_7)*signed(FMAP_19_31);
			MULT_32(18)<=signed(DIN_32_7)*signed(FMAP_19_32);
			MULT_33(18)<=signed(DIN_33_7)*signed(FMAP_19_33);
			MULT_34(18)<=signed(DIN_34_7)*signed(FMAP_19_34);
			MULT_35(18)<=signed(DIN_35_7)*signed(FMAP_19_35);
			MULT_36(18)<=signed(DIN_36_7)*signed(FMAP_19_36);
			MULT_37(18)<=signed(DIN_37_7)*signed(FMAP_19_37);
			MULT_38(18)<=signed(DIN_38_7)*signed(FMAP_19_38);
			MULT_39(18)<=signed(DIN_39_7)*signed(FMAP_19_39);
			MULT_40(18)<=signed(DIN_40_7)*signed(FMAP_19_40);
			MULT_41(18)<=signed(DIN_41_7)*signed(FMAP_19_41);
			MULT_42(18)<=signed(DIN_42_7)*signed(FMAP_19_42);
			MULT_43(18)<=signed(DIN_43_7)*signed(FMAP_19_43);
			MULT_44(18)<=signed(DIN_44_7)*signed(FMAP_19_44);
			MULT_45(18)<=signed(DIN_45_7)*signed(FMAP_19_45);
			MULT_46(18)<=signed(DIN_46_7)*signed(FMAP_19_46);
			MULT_47(18)<=signed(DIN_47_7)*signed(FMAP_19_47);
			MULT_48(18)<=signed(DIN_48_7)*signed(FMAP_19_48);
			MULT_49(18)<=signed(DIN_49_7)*signed(FMAP_19_49);
			MULT_50(18)<=signed(DIN_50_7)*signed(FMAP_19_50);
			MULT_51(18)<=signed(DIN_51_7)*signed(FMAP_19_51);
			MULT_52(18)<=signed(DIN_52_7)*signed(FMAP_19_52);
			MULT_53(18)<=signed(DIN_53_7)*signed(FMAP_19_53);
			MULT_54(18)<=signed(DIN_54_7)*signed(FMAP_19_54);
			MULT_55(18)<=signed(DIN_55_7)*signed(FMAP_19_55);
			MULT_56(18)<=signed(DIN_56_7)*signed(FMAP_19_56);
			MULT_57(18)<=signed(DIN_57_7)*signed(FMAP_19_57);
			MULT_58(18)<=signed(DIN_58_7)*signed(FMAP_19_58);
			MULT_59(18)<=signed(DIN_59_7)*signed(FMAP_19_59);
			MULT_60(18)<=signed(DIN_60_7)*signed(FMAP_19_60);
			MULT_61(18)<=signed(DIN_61_7)*signed(FMAP_19_61);
			MULT_62(18)<=signed(DIN_62_7)*signed(FMAP_19_62);
			MULT_63(18)<=signed(DIN_63_7)*signed(FMAP_19_63);
			MULT_64(18)<=signed(DIN_64_7)*signed(FMAP_19_64);
			MULT_65(18)<=signed(DIN_65_7)*signed(FMAP_19_65);
			MULT_66(18)<=signed(DIN_66_7)*signed(FMAP_19_66);
			MULT_67(18)<=signed(DIN_67_7)*signed(FMAP_19_67);
			MULT_68(18)<=signed(DIN_68_7)*signed(FMAP_19_68);
			MULT_69(18)<=signed(DIN_69_7)*signed(FMAP_19_69);
			MULT_70(18)<=signed(DIN_70_7)*signed(FMAP_19_70);
			MULT_71(18)<=signed(DIN_71_7)*signed(FMAP_19_71);
			MULT_72(18)<=signed(DIN_72_7)*signed(FMAP_19_72);
			MULT_73(18)<=signed(DIN_73_7)*signed(FMAP_19_73);
			MULT_74(18)<=signed(DIN_74_7)*signed(FMAP_19_74);
			MULT_75(18)<=signed(DIN_75_7)*signed(FMAP_19_75);
			MULT_76(18)<=signed(DIN_76_7)*signed(FMAP_19_76);
			MULT_77(18)<=signed(DIN_77_7)*signed(FMAP_19_77);
			MULT_78(18)<=signed(DIN_78_7)*signed(FMAP_19_78);
			MULT_79(18)<=signed(DIN_79_7)*signed(FMAP_19_79);
			MULT_80(18)<=signed(DIN_80_7)*signed(FMAP_19_80);
			MULT_81(18)<=signed(DIN_81_7)*signed(FMAP_19_81);
			MULT_82(18)<=signed(DIN_82_7)*signed(FMAP_19_82);
			MULT_83(18)<=signed(DIN_83_7)*signed(FMAP_19_83);
			MULT_84(18)<=signed(DIN_84_7)*signed(FMAP_19_84);
			MULT_85(18)<=signed(DIN_85_7)*signed(FMAP_19_85);
			MULT_86(18)<=signed(DIN_86_7)*signed(FMAP_19_86);
			MULT_87(18)<=signed(DIN_87_7)*signed(FMAP_19_87);
			MULT_88(18)<=signed(DIN_88_7)*signed(FMAP_19_88);
			MULT_89(18)<=signed(DIN_89_7)*signed(FMAP_19_89);
			MULT_90(18)<=signed(DIN_90_7)*signed(FMAP_19_90);
			MULT_91(18)<=signed(DIN_91_7)*signed(FMAP_19_91);
			MULT_92(18)<=signed(DIN_92_7)*signed(FMAP_19_92);
			MULT_93(18)<=signed(DIN_93_7)*signed(FMAP_19_93);
			MULT_94(18)<=signed(DIN_94_7)*signed(FMAP_19_94);
			MULT_95(18)<=signed(DIN_95_7)*signed(FMAP_19_95);
			MULT_96(18)<=signed(DIN_96_7)*signed(FMAP_19_96);
			MULT_97(18)<=signed(DIN_97_7)*signed(FMAP_19_97);
			MULT_98(18)<=signed(DIN_98_7)*signed(FMAP_19_98);
			MULT_99(18)<=signed(DIN_99_7)*signed(FMAP_19_99);
			MULT_100(18)<=signed(DIN_100_7)*signed(FMAP_19_100);
			MULT_101(18)<=signed(DIN_101_7)*signed(FMAP_19_101);
			MULT_102(18)<=signed(DIN_102_7)*signed(FMAP_19_102);
			MULT_103(18)<=signed(DIN_103_7)*signed(FMAP_19_103);
			MULT_104(18)<=signed(DIN_104_7)*signed(FMAP_19_104);
			MULT_105(18)<=signed(DIN_105_7)*signed(FMAP_19_105);
			MULT_106(18)<=signed(DIN_106_7)*signed(FMAP_19_106);
			MULT_107(18)<=signed(DIN_107_7)*signed(FMAP_19_107);
			MULT_108(18)<=signed(DIN_108_7)*signed(FMAP_19_108);
			MULT_109(18)<=signed(DIN_109_7)*signed(FMAP_19_109);
			MULT_110(18)<=signed(DIN_110_7)*signed(FMAP_19_110);
			MULT_111(18)<=signed(DIN_111_7)*signed(FMAP_19_111);
			MULT_112(18)<=signed(DIN_112_7)*signed(FMAP_19_112);
			MULT_113(18)<=signed(DIN_113_7)*signed(FMAP_19_113);
			MULT_114(18)<=signed(DIN_114_7)*signed(FMAP_19_114);
			MULT_115(18)<=signed(DIN_115_7)*signed(FMAP_19_115);
			MULT_116(18)<=signed(DIN_116_7)*signed(FMAP_19_116);
			MULT_117(18)<=signed(DIN_117_7)*signed(FMAP_19_117);
			MULT_118(18)<=signed(DIN_118_7)*signed(FMAP_19_118);
			MULT_119(18)<=signed(DIN_119_7)*signed(FMAP_19_119);
			MULT_120(18)<=signed(DIN_120_7)*signed(FMAP_19_120);

			MULT_1(19)<=signed(DIN_1_7)*signed(FMAP_20_1);
			MULT_2(19)<=signed(DIN_2_7)*signed(FMAP_20_2);
			MULT_3(19)<=signed(DIN_3_7)*signed(FMAP_20_3);
			MULT_4(19)<=signed(DIN_4_7)*signed(FMAP_20_4);
			MULT_5(19)<=signed(DIN_5_7)*signed(FMAP_20_5);
			MULT_6(19)<=signed(DIN_6_7)*signed(FMAP_20_6);
			MULT_7(19)<=signed(DIN_7_7)*signed(FMAP_20_7);
			MULT_8(19)<=signed(DIN_8_7)*signed(FMAP_20_8);
			MULT_9(19)<=signed(DIN_9_7)*signed(FMAP_20_9);
			MULT_10(19)<=signed(DIN_10_7)*signed(FMAP_20_10);
			MULT_11(19)<=signed(DIN_11_7)*signed(FMAP_20_11);
			MULT_12(19)<=signed(DIN_12_7)*signed(FMAP_20_12);
			MULT_13(19)<=signed(DIN_13_7)*signed(FMAP_20_13);
			MULT_14(19)<=signed(DIN_14_7)*signed(FMAP_20_14);
			MULT_15(19)<=signed(DIN_15_7)*signed(FMAP_20_15);
			MULT_16(19)<=signed(DIN_16_7)*signed(FMAP_20_16);
			MULT_17(19)<=signed(DIN_17_7)*signed(FMAP_20_17);
			MULT_18(19)<=signed(DIN_18_7)*signed(FMAP_20_18);
			MULT_19(19)<=signed(DIN_19_7)*signed(FMAP_20_19);
			MULT_20(19)<=signed(DIN_20_7)*signed(FMAP_20_20);
			MULT_21(19)<=signed(DIN_21_7)*signed(FMAP_20_21);
			MULT_22(19)<=signed(DIN_22_7)*signed(FMAP_20_22);
			MULT_23(19)<=signed(DIN_23_7)*signed(FMAP_20_23);
			MULT_24(19)<=signed(DIN_24_7)*signed(FMAP_20_24);
			MULT_25(19)<=signed(DIN_25_7)*signed(FMAP_20_25);
			MULT_26(19)<=signed(DIN_26_7)*signed(FMAP_20_26);
			MULT_27(19)<=signed(DIN_27_7)*signed(FMAP_20_27);
			MULT_28(19)<=signed(DIN_28_7)*signed(FMAP_20_28);
			MULT_29(19)<=signed(DIN_29_7)*signed(FMAP_20_29);
			MULT_30(19)<=signed(DIN_30_7)*signed(FMAP_20_30);
			MULT_31(19)<=signed(DIN_31_7)*signed(FMAP_20_31);
			MULT_32(19)<=signed(DIN_32_7)*signed(FMAP_20_32);
			MULT_33(19)<=signed(DIN_33_7)*signed(FMAP_20_33);
			MULT_34(19)<=signed(DIN_34_7)*signed(FMAP_20_34);
			MULT_35(19)<=signed(DIN_35_7)*signed(FMAP_20_35);
			MULT_36(19)<=signed(DIN_36_7)*signed(FMAP_20_36);
			MULT_37(19)<=signed(DIN_37_7)*signed(FMAP_20_37);
			MULT_38(19)<=signed(DIN_38_7)*signed(FMAP_20_38);
			MULT_39(19)<=signed(DIN_39_7)*signed(FMAP_20_39);
			MULT_40(19)<=signed(DIN_40_7)*signed(FMAP_20_40);
			MULT_41(19)<=signed(DIN_41_7)*signed(FMAP_20_41);
			MULT_42(19)<=signed(DIN_42_7)*signed(FMAP_20_42);
			MULT_43(19)<=signed(DIN_43_7)*signed(FMAP_20_43);
			MULT_44(19)<=signed(DIN_44_7)*signed(FMAP_20_44);
			MULT_45(19)<=signed(DIN_45_7)*signed(FMAP_20_45);
			MULT_46(19)<=signed(DIN_46_7)*signed(FMAP_20_46);
			MULT_47(19)<=signed(DIN_47_7)*signed(FMAP_20_47);
			MULT_48(19)<=signed(DIN_48_7)*signed(FMAP_20_48);
			MULT_49(19)<=signed(DIN_49_7)*signed(FMAP_20_49);
			MULT_50(19)<=signed(DIN_50_7)*signed(FMAP_20_50);
			MULT_51(19)<=signed(DIN_51_7)*signed(FMAP_20_51);
			MULT_52(19)<=signed(DIN_52_7)*signed(FMAP_20_52);
			MULT_53(19)<=signed(DIN_53_7)*signed(FMAP_20_53);
			MULT_54(19)<=signed(DIN_54_7)*signed(FMAP_20_54);
			MULT_55(19)<=signed(DIN_55_7)*signed(FMAP_20_55);
			MULT_56(19)<=signed(DIN_56_7)*signed(FMAP_20_56);
			MULT_57(19)<=signed(DIN_57_7)*signed(FMAP_20_57);
			MULT_58(19)<=signed(DIN_58_7)*signed(FMAP_20_58);
			MULT_59(19)<=signed(DIN_59_7)*signed(FMAP_20_59);
			MULT_60(19)<=signed(DIN_60_7)*signed(FMAP_20_60);
			MULT_61(19)<=signed(DIN_61_7)*signed(FMAP_20_61);
			MULT_62(19)<=signed(DIN_62_7)*signed(FMAP_20_62);
			MULT_63(19)<=signed(DIN_63_7)*signed(FMAP_20_63);
			MULT_64(19)<=signed(DIN_64_7)*signed(FMAP_20_64);
			MULT_65(19)<=signed(DIN_65_7)*signed(FMAP_20_65);
			MULT_66(19)<=signed(DIN_66_7)*signed(FMAP_20_66);
			MULT_67(19)<=signed(DIN_67_7)*signed(FMAP_20_67);
			MULT_68(19)<=signed(DIN_68_7)*signed(FMAP_20_68);
			MULT_69(19)<=signed(DIN_69_7)*signed(FMAP_20_69);
			MULT_70(19)<=signed(DIN_70_7)*signed(FMAP_20_70);
			MULT_71(19)<=signed(DIN_71_7)*signed(FMAP_20_71);
			MULT_72(19)<=signed(DIN_72_7)*signed(FMAP_20_72);
			MULT_73(19)<=signed(DIN_73_7)*signed(FMAP_20_73);
			MULT_74(19)<=signed(DIN_74_7)*signed(FMAP_20_74);
			MULT_75(19)<=signed(DIN_75_7)*signed(FMAP_20_75);
			MULT_76(19)<=signed(DIN_76_7)*signed(FMAP_20_76);
			MULT_77(19)<=signed(DIN_77_7)*signed(FMAP_20_77);
			MULT_78(19)<=signed(DIN_78_7)*signed(FMAP_20_78);
			MULT_79(19)<=signed(DIN_79_7)*signed(FMAP_20_79);
			MULT_80(19)<=signed(DIN_80_7)*signed(FMAP_20_80);
			MULT_81(19)<=signed(DIN_81_7)*signed(FMAP_20_81);
			MULT_82(19)<=signed(DIN_82_7)*signed(FMAP_20_82);
			MULT_83(19)<=signed(DIN_83_7)*signed(FMAP_20_83);
			MULT_84(19)<=signed(DIN_84_7)*signed(FMAP_20_84);
			MULT_85(19)<=signed(DIN_85_7)*signed(FMAP_20_85);
			MULT_86(19)<=signed(DIN_86_7)*signed(FMAP_20_86);
			MULT_87(19)<=signed(DIN_87_7)*signed(FMAP_20_87);
			MULT_88(19)<=signed(DIN_88_7)*signed(FMAP_20_88);
			MULT_89(19)<=signed(DIN_89_7)*signed(FMAP_20_89);
			MULT_90(19)<=signed(DIN_90_7)*signed(FMAP_20_90);
			MULT_91(19)<=signed(DIN_91_7)*signed(FMAP_20_91);
			MULT_92(19)<=signed(DIN_92_7)*signed(FMAP_20_92);
			MULT_93(19)<=signed(DIN_93_7)*signed(FMAP_20_93);
			MULT_94(19)<=signed(DIN_94_7)*signed(FMAP_20_94);
			MULT_95(19)<=signed(DIN_95_7)*signed(FMAP_20_95);
			MULT_96(19)<=signed(DIN_96_7)*signed(FMAP_20_96);
			MULT_97(19)<=signed(DIN_97_7)*signed(FMAP_20_97);
			MULT_98(19)<=signed(DIN_98_7)*signed(FMAP_20_98);
			MULT_99(19)<=signed(DIN_99_7)*signed(FMAP_20_99);
			MULT_100(19)<=signed(DIN_100_7)*signed(FMAP_20_100);
			MULT_101(19)<=signed(DIN_101_7)*signed(FMAP_20_101);
			MULT_102(19)<=signed(DIN_102_7)*signed(FMAP_20_102);
			MULT_103(19)<=signed(DIN_103_7)*signed(FMAP_20_103);
			MULT_104(19)<=signed(DIN_104_7)*signed(FMAP_20_104);
			MULT_105(19)<=signed(DIN_105_7)*signed(FMAP_20_105);
			MULT_106(19)<=signed(DIN_106_7)*signed(FMAP_20_106);
			MULT_107(19)<=signed(DIN_107_7)*signed(FMAP_20_107);
			MULT_108(19)<=signed(DIN_108_7)*signed(FMAP_20_108);
			MULT_109(19)<=signed(DIN_109_7)*signed(FMAP_20_109);
			MULT_110(19)<=signed(DIN_110_7)*signed(FMAP_20_110);
			MULT_111(19)<=signed(DIN_111_7)*signed(FMAP_20_111);
			MULT_112(19)<=signed(DIN_112_7)*signed(FMAP_20_112);
			MULT_113(19)<=signed(DIN_113_7)*signed(FMAP_20_113);
			MULT_114(19)<=signed(DIN_114_7)*signed(FMAP_20_114);
			MULT_115(19)<=signed(DIN_115_7)*signed(FMAP_20_115);
			MULT_116(19)<=signed(DIN_116_7)*signed(FMAP_20_116);
			MULT_117(19)<=signed(DIN_117_7)*signed(FMAP_20_117);
			MULT_118(19)<=signed(DIN_118_7)*signed(FMAP_20_118);
			MULT_119(19)<=signed(DIN_119_7)*signed(FMAP_20_119);
			MULT_120(19)<=signed(DIN_120_7)*signed(FMAP_20_120);

			MULT_1(20)<=signed(DIN_1_7)*signed(FMAP_21_1);
			MULT_2(20)<=signed(DIN_2_7)*signed(FMAP_21_2);
			MULT_3(20)<=signed(DIN_3_7)*signed(FMAP_21_3);
			MULT_4(20)<=signed(DIN_4_7)*signed(FMAP_21_4);
			MULT_5(20)<=signed(DIN_5_7)*signed(FMAP_21_5);
			MULT_6(20)<=signed(DIN_6_7)*signed(FMAP_21_6);
			MULT_7(20)<=signed(DIN_7_7)*signed(FMAP_21_7);
			MULT_8(20)<=signed(DIN_8_7)*signed(FMAP_21_8);
			MULT_9(20)<=signed(DIN_9_7)*signed(FMAP_21_9);
			MULT_10(20)<=signed(DIN_10_7)*signed(FMAP_21_10);
			MULT_11(20)<=signed(DIN_11_7)*signed(FMAP_21_11);
			MULT_12(20)<=signed(DIN_12_7)*signed(FMAP_21_12);
			MULT_13(20)<=signed(DIN_13_7)*signed(FMAP_21_13);
			MULT_14(20)<=signed(DIN_14_7)*signed(FMAP_21_14);
			MULT_15(20)<=signed(DIN_15_7)*signed(FMAP_21_15);
			MULT_16(20)<=signed(DIN_16_7)*signed(FMAP_21_16);
			MULT_17(20)<=signed(DIN_17_7)*signed(FMAP_21_17);
			MULT_18(20)<=signed(DIN_18_7)*signed(FMAP_21_18);
			MULT_19(20)<=signed(DIN_19_7)*signed(FMAP_21_19);
			MULT_20(20)<=signed(DIN_20_7)*signed(FMAP_21_20);
			MULT_21(20)<=signed(DIN_21_7)*signed(FMAP_21_21);
			MULT_22(20)<=signed(DIN_22_7)*signed(FMAP_21_22);
			MULT_23(20)<=signed(DIN_23_7)*signed(FMAP_21_23);
			MULT_24(20)<=signed(DIN_24_7)*signed(FMAP_21_24);
			MULT_25(20)<=signed(DIN_25_7)*signed(FMAP_21_25);
			MULT_26(20)<=signed(DIN_26_7)*signed(FMAP_21_26);
			MULT_27(20)<=signed(DIN_27_7)*signed(FMAP_21_27);
			MULT_28(20)<=signed(DIN_28_7)*signed(FMAP_21_28);
			MULT_29(20)<=signed(DIN_29_7)*signed(FMAP_21_29);
			MULT_30(20)<=signed(DIN_30_7)*signed(FMAP_21_30);
			MULT_31(20)<=signed(DIN_31_7)*signed(FMAP_21_31);
			MULT_32(20)<=signed(DIN_32_7)*signed(FMAP_21_32);
			MULT_33(20)<=signed(DIN_33_7)*signed(FMAP_21_33);
			MULT_34(20)<=signed(DIN_34_7)*signed(FMAP_21_34);
			MULT_35(20)<=signed(DIN_35_7)*signed(FMAP_21_35);
			MULT_36(20)<=signed(DIN_36_7)*signed(FMAP_21_36);
			MULT_37(20)<=signed(DIN_37_7)*signed(FMAP_21_37);
			MULT_38(20)<=signed(DIN_38_7)*signed(FMAP_21_38);
			MULT_39(20)<=signed(DIN_39_7)*signed(FMAP_21_39);
			MULT_40(20)<=signed(DIN_40_7)*signed(FMAP_21_40);
			MULT_41(20)<=signed(DIN_41_7)*signed(FMAP_21_41);
			MULT_42(20)<=signed(DIN_42_7)*signed(FMAP_21_42);
			MULT_43(20)<=signed(DIN_43_7)*signed(FMAP_21_43);
			MULT_44(20)<=signed(DIN_44_7)*signed(FMAP_21_44);
			MULT_45(20)<=signed(DIN_45_7)*signed(FMAP_21_45);
			MULT_46(20)<=signed(DIN_46_7)*signed(FMAP_21_46);
			MULT_47(20)<=signed(DIN_47_7)*signed(FMAP_21_47);
			MULT_48(20)<=signed(DIN_48_7)*signed(FMAP_21_48);
			MULT_49(20)<=signed(DIN_49_7)*signed(FMAP_21_49);
			MULT_50(20)<=signed(DIN_50_7)*signed(FMAP_21_50);
			MULT_51(20)<=signed(DIN_51_7)*signed(FMAP_21_51);
			MULT_52(20)<=signed(DIN_52_7)*signed(FMAP_21_52);
			MULT_53(20)<=signed(DIN_53_7)*signed(FMAP_21_53);
			MULT_54(20)<=signed(DIN_54_7)*signed(FMAP_21_54);
			MULT_55(20)<=signed(DIN_55_7)*signed(FMAP_21_55);
			MULT_56(20)<=signed(DIN_56_7)*signed(FMAP_21_56);
			MULT_57(20)<=signed(DIN_57_7)*signed(FMAP_21_57);
			MULT_58(20)<=signed(DIN_58_7)*signed(FMAP_21_58);
			MULT_59(20)<=signed(DIN_59_7)*signed(FMAP_21_59);
			MULT_60(20)<=signed(DIN_60_7)*signed(FMAP_21_60);
			MULT_61(20)<=signed(DIN_61_7)*signed(FMAP_21_61);
			MULT_62(20)<=signed(DIN_62_7)*signed(FMAP_21_62);
			MULT_63(20)<=signed(DIN_63_7)*signed(FMAP_21_63);
			MULT_64(20)<=signed(DIN_64_7)*signed(FMAP_21_64);
			MULT_65(20)<=signed(DIN_65_7)*signed(FMAP_21_65);
			MULT_66(20)<=signed(DIN_66_7)*signed(FMAP_21_66);
			MULT_67(20)<=signed(DIN_67_7)*signed(FMAP_21_67);
			MULT_68(20)<=signed(DIN_68_7)*signed(FMAP_21_68);
			MULT_69(20)<=signed(DIN_69_7)*signed(FMAP_21_69);
			MULT_70(20)<=signed(DIN_70_7)*signed(FMAP_21_70);
			MULT_71(20)<=signed(DIN_71_7)*signed(FMAP_21_71);
			MULT_72(20)<=signed(DIN_72_7)*signed(FMAP_21_72);
			MULT_73(20)<=signed(DIN_73_7)*signed(FMAP_21_73);
			MULT_74(20)<=signed(DIN_74_7)*signed(FMAP_21_74);
			MULT_75(20)<=signed(DIN_75_7)*signed(FMAP_21_75);
			MULT_76(20)<=signed(DIN_76_7)*signed(FMAP_21_76);
			MULT_77(20)<=signed(DIN_77_7)*signed(FMAP_21_77);
			MULT_78(20)<=signed(DIN_78_7)*signed(FMAP_21_78);
			MULT_79(20)<=signed(DIN_79_7)*signed(FMAP_21_79);
			MULT_80(20)<=signed(DIN_80_7)*signed(FMAP_21_80);
			MULT_81(20)<=signed(DIN_81_7)*signed(FMAP_21_81);
			MULT_82(20)<=signed(DIN_82_7)*signed(FMAP_21_82);
			MULT_83(20)<=signed(DIN_83_7)*signed(FMAP_21_83);
			MULT_84(20)<=signed(DIN_84_7)*signed(FMAP_21_84);
			MULT_85(20)<=signed(DIN_85_7)*signed(FMAP_21_85);
			MULT_86(20)<=signed(DIN_86_7)*signed(FMAP_21_86);
			MULT_87(20)<=signed(DIN_87_7)*signed(FMAP_21_87);
			MULT_88(20)<=signed(DIN_88_7)*signed(FMAP_21_88);
			MULT_89(20)<=signed(DIN_89_7)*signed(FMAP_21_89);
			MULT_90(20)<=signed(DIN_90_7)*signed(FMAP_21_90);
			MULT_91(20)<=signed(DIN_91_7)*signed(FMAP_21_91);
			MULT_92(20)<=signed(DIN_92_7)*signed(FMAP_21_92);
			MULT_93(20)<=signed(DIN_93_7)*signed(FMAP_21_93);
			MULT_94(20)<=signed(DIN_94_7)*signed(FMAP_21_94);
			MULT_95(20)<=signed(DIN_95_7)*signed(FMAP_21_95);
			MULT_96(20)<=signed(DIN_96_7)*signed(FMAP_21_96);
			MULT_97(20)<=signed(DIN_97_7)*signed(FMAP_21_97);
			MULT_98(20)<=signed(DIN_98_7)*signed(FMAP_21_98);
			MULT_99(20)<=signed(DIN_99_7)*signed(FMAP_21_99);
			MULT_100(20)<=signed(DIN_100_7)*signed(FMAP_21_100);
			MULT_101(20)<=signed(DIN_101_7)*signed(FMAP_21_101);
			MULT_102(20)<=signed(DIN_102_7)*signed(FMAP_21_102);
			MULT_103(20)<=signed(DIN_103_7)*signed(FMAP_21_103);
			MULT_104(20)<=signed(DIN_104_7)*signed(FMAP_21_104);
			MULT_105(20)<=signed(DIN_105_7)*signed(FMAP_21_105);
			MULT_106(20)<=signed(DIN_106_7)*signed(FMAP_21_106);
			MULT_107(20)<=signed(DIN_107_7)*signed(FMAP_21_107);
			MULT_108(20)<=signed(DIN_108_7)*signed(FMAP_21_108);
			MULT_109(20)<=signed(DIN_109_7)*signed(FMAP_21_109);
			MULT_110(20)<=signed(DIN_110_7)*signed(FMAP_21_110);
			MULT_111(20)<=signed(DIN_111_7)*signed(FMAP_21_111);
			MULT_112(20)<=signed(DIN_112_7)*signed(FMAP_21_112);
			MULT_113(20)<=signed(DIN_113_7)*signed(FMAP_21_113);
			MULT_114(20)<=signed(DIN_114_7)*signed(FMAP_21_114);
			MULT_115(20)<=signed(DIN_115_7)*signed(FMAP_21_115);
			MULT_116(20)<=signed(DIN_116_7)*signed(FMAP_21_116);
			MULT_117(20)<=signed(DIN_117_7)*signed(FMAP_21_117);
			MULT_118(20)<=signed(DIN_118_7)*signed(FMAP_21_118);
			MULT_119(20)<=signed(DIN_119_7)*signed(FMAP_21_119);
			MULT_120(20)<=signed(DIN_120_7)*signed(FMAP_21_120);

			MULT_1(21)<=signed(DIN_1_7)*signed(FMAP_22_1);
			MULT_2(21)<=signed(DIN_2_7)*signed(FMAP_22_2);
			MULT_3(21)<=signed(DIN_3_7)*signed(FMAP_22_3);
			MULT_4(21)<=signed(DIN_4_7)*signed(FMAP_22_4);
			MULT_5(21)<=signed(DIN_5_7)*signed(FMAP_22_5);
			MULT_6(21)<=signed(DIN_6_7)*signed(FMAP_22_6);
			MULT_7(21)<=signed(DIN_7_7)*signed(FMAP_22_7);
			MULT_8(21)<=signed(DIN_8_7)*signed(FMAP_22_8);
			MULT_9(21)<=signed(DIN_9_7)*signed(FMAP_22_9);
			MULT_10(21)<=signed(DIN_10_7)*signed(FMAP_22_10);
			MULT_11(21)<=signed(DIN_11_7)*signed(FMAP_22_11);
			MULT_12(21)<=signed(DIN_12_7)*signed(FMAP_22_12);
			MULT_13(21)<=signed(DIN_13_7)*signed(FMAP_22_13);
			MULT_14(21)<=signed(DIN_14_7)*signed(FMAP_22_14);
			MULT_15(21)<=signed(DIN_15_7)*signed(FMAP_22_15);
			MULT_16(21)<=signed(DIN_16_7)*signed(FMAP_22_16);
			MULT_17(21)<=signed(DIN_17_7)*signed(FMAP_22_17);
			MULT_18(21)<=signed(DIN_18_7)*signed(FMAP_22_18);
			MULT_19(21)<=signed(DIN_19_7)*signed(FMAP_22_19);
			MULT_20(21)<=signed(DIN_20_7)*signed(FMAP_22_20);
			MULT_21(21)<=signed(DIN_21_7)*signed(FMAP_22_21);
			MULT_22(21)<=signed(DIN_22_7)*signed(FMAP_22_22);
			MULT_23(21)<=signed(DIN_23_7)*signed(FMAP_22_23);
			MULT_24(21)<=signed(DIN_24_7)*signed(FMAP_22_24);
			MULT_25(21)<=signed(DIN_25_7)*signed(FMAP_22_25);
			MULT_26(21)<=signed(DIN_26_7)*signed(FMAP_22_26);
			MULT_27(21)<=signed(DIN_27_7)*signed(FMAP_22_27);
			MULT_28(21)<=signed(DIN_28_7)*signed(FMAP_22_28);
			MULT_29(21)<=signed(DIN_29_7)*signed(FMAP_22_29);
			MULT_30(21)<=signed(DIN_30_7)*signed(FMAP_22_30);
			MULT_31(21)<=signed(DIN_31_7)*signed(FMAP_22_31);
			MULT_32(21)<=signed(DIN_32_7)*signed(FMAP_22_32);
			MULT_33(21)<=signed(DIN_33_7)*signed(FMAP_22_33);
			MULT_34(21)<=signed(DIN_34_7)*signed(FMAP_22_34);
			MULT_35(21)<=signed(DIN_35_7)*signed(FMAP_22_35);
			MULT_36(21)<=signed(DIN_36_7)*signed(FMAP_22_36);
			MULT_37(21)<=signed(DIN_37_7)*signed(FMAP_22_37);
			MULT_38(21)<=signed(DIN_38_7)*signed(FMAP_22_38);
			MULT_39(21)<=signed(DIN_39_7)*signed(FMAP_22_39);
			MULT_40(21)<=signed(DIN_40_7)*signed(FMAP_22_40);
			MULT_41(21)<=signed(DIN_41_7)*signed(FMAP_22_41);
			MULT_42(21)<=signed(DIN_42_7)*signed(FMAP_22_42);
			MULT_43(21)<=signed(DIN_43_7)*signed(FMAP_22_43);
			MULT_44(21)<=signed(DIN_44_7)*signed(FMAP_22_44);
			MULT_45(21)<=signed(DIN_45_7)*signed(FMAP_22_45);
			MULT_46(21)<=signed(DIN_46_7)*signed(FMAP_22_46);
			MULT_47(21)<=signed(DIN_47_7)*signed(FMAP_22_47);
			MULT_48(21)<=signed(DIN_48_7)*signed(FMAP_22_48);
			MULT_49(21)<=signed(DIN_49_7)*signed(FMAP_22_49);
			MULT_50(21)<=signed(DIN_50_7)*signed(FMAP_22_50);
			MULT_51(21)<=signed(DIN_51_7)*signed(FMAP_22_51);
			MULT_52(21)<=signed(DIN_52_7)*signed(FMAP_22_52);
			MULT_53(21)<=signed(DIN_53_7)*signed(FMAP_22_53);
			MULT_54(21)<=signed(DIN_54_7)*signed(FMAP_22_54);
			MULT_55(21)<=signed(DIN_55_7)*signed(FMAP_22_55);
			MULT_56(21)<=signed(DIN_56_7)*signed(FMAP_22_56);
			MULT_57(21)<=signed(DIN_57_7)*signed(FMAP_22_57);
			MULT_58(21)<=signed(DIN_58_7)*signed(FMAP_22_58);
			MULT_59(21)<=signed(DIN_59_7)*signed(FMAP_22_59);
			MULT_60(21)<=signed(DIN_60_7)*signed(FMAP_22_60);
			MULT_61(21)<=signed(DIN_61_7)*signed(FMAP_22_61);
			MULT_62(21)<=signed(DIN_62_7)*signed(FMAP_22_62);
			MULT_63(21)<=signed(DIN_63_7)*signed(FMAP_22_63);
			MULT_64(21)<=signed(DIN_64_7)*signed(FMAP_22_64);
			MULT_65(21)<=signed(DIN_65_7)*signed(FMAP_22_65);
			MULT_66(21)<=signed(DIN_66_7)*signed(FMAP_22_66);
			MULT_67(21)<=signed(DIN_67_7)*signed(FMAP_22_67);
			MULT_68(21)<=signed(DIN_68_7)*signed(FMAP_22_68);
			MULT_69(21)<=signed(DIN_69_7)*signed(FMAP_22_69);
			MULT_70(21)<=signed(DIN_70_7)*signed(FMAP_22_70);
			MULT_71(21)<=signed(DIN_71_7)*signed(FMAP_22_71);
			MULT_72(21)<=signed(DIN_72_7)*signed(FMAP_22_72);
			MULT_73(21)<=signed(DIN_73_7)*signed(FMAP_22_73);
			MULT_74(21)<=signed(DIN_74_7)*signed(FMAP_22_74);
			MULT_75(21)<=signed(DIN_75_7)*signed(FMAP_22_75);
			MULT_76(21)<=signed(DIN_76_7)*signed(FMAP_22_76);
			MULT_77(21)<=signed(DIN_77_7)*signed(FMAP_22_77);
			MULT_78(21)<=signed(DIN_78_7)*signed(FMAP_22_78);
			MULT_79(21)<=signed(DIN_79_7)*signed(FMAP_22_79);
			MULT_80(21)<=signed(DIN_80_7)*signed(FMAP_22_80);
			MULT_81(21)<=signed(DIN_81_7)*signed(FMAP_22_81);
			MULT_82(21)<=signed(DIN_82_7)*signed(FMAP_22_82);
			MULT_83(21)<=signed(DIN_83_7)*signed(FMAP_22_83);
			MULT_84(21)<=signed(DIN_84_7)*signed(FMAP_22_84);
			MULT_85(21)<=signed(DIN_85_7)*signed(FMAP_22_85);
			MULT_86(21)<=signed(DIN_86_7)*signed(FMAP_22_86);
			MULT_87(21)<=signed(DIN_87_7)*signed(FMAP_22_87);
			MULT_88(21)<=signed(DIN_88_7)*signed(FMAP_22_88);
			MULT_89(21)<=signed(DIN_89_7)*signed(FMAP_22_89);
			MULT_90(21)<=signed(DIN_90_7)*signed(FMAP_22_90);
			MULT_91(21)<=signed(DIN_91_7)*signed(FMAP_22_91);
			MULT_92(21)<=signed(DIN_92_7)*signed(FMAP_22_92);
			MULT_93(21)<=signed(DIN_93_7)*signed(FMAP_22_93);
			MULT_94(21)<=signed(DIN_94_7)*signed(FMAP_22_94);
			MULT_95(21)<=signed(DIN_95_7)*signed(FMAP_22_95);
			MULT_96(21)<=signed(DIN_96_7)*signed(FMAP_22_96);
			MULT_97(21)<=signed(DIN_97_7)*signed(FMAP_22_97);
			MULT_98(21)<=signed(DIN_98_7)*signed(FMAP_22_98);
			MULT_99(21)<=signed(DIN_99_7)*signed(FMAP_22_99);
			MULT_100(21)<=signed(DIN_100_7)*signed(FMAP_22_100);
			MULT_101(21)<=signed(DIN_101_7)*signed(FMAP_22_101);
			MULT_102(21)<=signed(DIN_102_7)*signed(FMAP_22_102);
			MULT_103(21)<=signed(DIN_103_7)*signed(FMAP_22_103);
			MULT_104(21)<=signed(DIN_104_7)*signed(FMAP_22_104);
			MULT_105(21)<=signed(DIN_105_7)*signed(FMAP_22_105);
			MULT_106(21)<=signed(DIN_106_7)*signed(FMAP_22_106);
			MULT_107(21)<=signed(DIN_107_7)*signed(FMAP_22_107);
			MULT_108(21)<=signed(DIN_108_7)*signed(FMAP_22_108);
			MULT_109(21)<=signed(DIN_109_7)*signed(FMAP_22_109);
			MULT_110(21)<=signed(DIN_110_7)*signed(FMAP_22_110);
			MULT_111(21)<=signed(DIN_111_7)*signed(FMAP_22_111);
			MULT_112(21)<=signed(DIN_112_7)*signed(FMAP_22_112);
			MULT_113(21)<=signed(DIN_113_7)*signed(FMAP_22_113);
			MULT_114(21)<=signed(DIN_114_7)*signed(FMAP_22_114);
			MULT_115(21)<=signed(DIN_115_7)*signed(FMAP_22_115);
			MULT_116(21)<=signed(DIN_116_7)*signed(FMAP_22_116);
			MULT_117(21)<=signed(DIN_117_7)*signed(FMAP_22_117);
			MULT_118(21)<=signed(DIN_118_7)*signed(FMAP_22_118);
			MULT_119(21)<=signed(DIN_119_7)*signed(FMAP_22_119);
			MULT_120(21)<=signed(DIN_120_7)*signed(FMAP_22_120);

			MULT_1(22)<=signed(DIN_1_7)*signed(FMAP_23_1);
			MULT_2(22)<=signed(DIN_2_7)*signed(FMAP_23_2);
			MULT_3(22)<=signed(DIN_3_7)*signed(FMAP_23_3);
			MULT_4(22)<=signed(DIN_4_7)*signed(FMAP_23_4);
			MULT_5(22)<=signed(DIN_5_7)*signed(FMAP_23_5);
			MULT_6(22)<=signed(DIN_6_7)*signed(FMAP_23_6);
			MULT_7(22)<=signed(DIN_7_7)*signed(FMAP_23_7);
			MULT_8(22)<=signed(DIN_8_7)*signed(FMAP_23_8);
			MULT_9(22)<=signed(DIN_9_7)*signed(FMAP_23_9);
			MULT_10(22)<=signed(DIN_10_7)*signed(FMAP_23_10);
			MULT_11(22)<=signed(DIN_11_7)*signed(FMAP_23_11);
			MULT_12(22)<=signed(DIN_12_7)*signed(FMAP_23_12);
			MULT_13(22)<=signed(DIN_13_7)*signed(FMAP_23_13);
			MULT_14(22)<=signed(DIN_14_7)*signed(FMAP_23_14);
			MULT_15(22)<=signed(DIN_15_7)*signed(FMAP_23_15);
			MULT_16(22)<=signed(DIN_16_7)*signed(FMAP_23_16);
			MULT_17(22)<=signed(DIN_17_7)*signed(FMAP_23_17);
			MULT_18(22)<=signed(DIN_18_7)*signed(FMAP_23_18);
			MULT_19(22)<=signed(DIN_19_7)*signed(FMAP_23_19);
			MULT_20(22)<=signed(DIN_20_7)*signed(FMAP_23_20);
			MULT_21(22)<=signed(DIN_21_7)*signed(FMAP_23_21);
			MULT_22(22)<=signed(DIN_22_7)*signed(FMAP_23_22);
			MULT_23(22)<=signed(DIN_23_7)*signed(FMAP_23_23);
			MULT_24(22)<=signed(DIN_24_7)*signed(FMAP_23_24);
			MULT_25(22)<=signed(DIN_25_7)*signed(FMAP_23_25);
			MULT_26(22)<=signed(DIN_26_7)*signed(FMAP_23_26);
			MULT_27(22)<=signed(DIN_27_7)*signed(FMAP_23_27);
			MULT_28(22)<=signed(DIN_28_7)*signed(FMAP_23_28);
			MULT_29(22)<=signed(DIN_29_7)*signed(FMAP_23_29);
			MULT_30(22)<=signed(DIN_30_7)*signed(FMAP_23_30);
			MULT_31(22)<=signed(DIN_31_7)*signed(FMAP_23_31);
			MULT_32(22)<=signed(DIN_32_7)*signed(FMAP_23_32);
			MULT_33(22)<=signed(DIN_33_7)*signed(FMAP_23_33);
			MULT_34(22)<=signed(DIN_34_7)*signed(FMAP_23_34);
			MULT_35(22)<=signed(DIN_35_7)*signed(FMAP_23_35);
			MULT_36(22)<=signed(DIN_36_7)*signed(FMAP_23_36);
			MULT_37(22)<=signed(DIN_37_7)*signed(FMAP_23_37);
			MULT_38(22)<=signed(DIN_38_7)*signed(FMAP_23_38);
			MULT_39(22)<=signed(DIN_39_7)*signed(FMAP_23_39);
			MULT_40(22)<=signed(DIN_40_7)*signed(FMAP_23_40);
			MULT_41(22)<=signed(DIN_41_7)*signed(FMAP_23_41);
			MULT_42(22)<=signed(DIN_42_7)*signed(FMAP_23_42);
			MULT_43(22)<=signed(DIN_43_7)*signed(FMAP_23_43);
			MULT_44(22)<=signed(DIN_44_7)*signed(FMAP_23_44);
			MULT_45(22)<=signed(DIN_45_7)*signed(FMAP_23_45);
			MULT_46(22)<=signed(DIN_46_7)*signed(FMAP_23_46);
			MULT_47(22)<=signed(DIN_47_7)*signed(FMAP_23_47);
			MULT_48(22)<=signed(DIN_48_7)*signed(FMAP_23_48);
			MULT_49(22)<=signed(DIN_49_7)*signed(FMAP_23_49);
			MULT_50(22)<=signed(DIN_50_7)*signed(FMAP_23_50);
			MULT_51(22)<=signed(DIN_51_7)*signed(FMAP_23_51);
			MULT_52(22)<=signed(DIN_52_7)*signed(FMAP_23_52);
			MULT_53(22)<=signed(DIN_53_7)*signed(FMAP_23_53);
			MULT_54(22)<=signed(DIN_54_7)*signed(FMAP_23_54);
			MULT_55(22)<=signed(DIN_55_7)*signed(FMAP_23_55);
			MULT_56(22)<=signed(DIN_56_7)*signed(FMAP_23_56);
			MULT_57(22)<=signed(DIN_57_7)*signed(FMAP_23_57);
			MULT_58(22)<=signed(DIN_58_7)*signed(FMAP_23_58);
			MULT_59(22)<=signed(DIN_59_7)*signed(FMAP_23_59);
			MULT_60(22)<=signed(DIN_60_7)*signed(FMAP_23_60);
			MULT_61(22)<=signed(DIN_61_7)*signed(FMAP_23_61);
			MULT_62(22)<=signed(DIN_62_7)*signed(FMAP_23_62);
			MULT_63(22)<=signed(DIN_63_7)*signed(FMAP_23_63);
			MULT_64(22)<=signed(DIN_64_7)*signed(FMAP_23_64);
			MULT_65(22)<=signed(DIN_65_7)*signed(FMAP_23_65);
			MULT_66(22)<=signed(DIN_66_7)*signed(FMAP_23_66);
			MULT_67(22)<=signed(DIN_67_7)*signed(FMAP_23_67);
			MULT_68(22)<=signed(DIN_68_7)*signed(FMAP_23_68);
			MULT_69(22)<=signed(DIN_69_7)*signed(FMAP_23_69);
			MULT_70(22)<=signed(DIN_70_7)*signed(FMAP_23_70);
			MULT_71(22)<=signed(DIN_71_7)*signed(FMAP_23_71);
			MULT_72(22)<=signed(DIN_72_7)*signed(FMAP_23_72);
			MULT_73(22)<=signed(DIN_73_7)*signed(FMAP_23_73);
			MULT_74(22)<=signed(DIN_74_7)*signed(FMAP_23_74);
			MULT_75(22)<=signed(DIN_75_7)*signed(FMAP_23_75);
			MULT_76(22)<=signed(DIN_76_7)*signed(FMAP_23_76);
			MULT_77(22)<=signed(DIN_77_7)*signed(FMAP_23_77);
			MULT_78(22)<=signed(DIN_78_7)*signed(FMAP_23_78);
			MULT_79(22)<=signed(DIN_79_7)*signed(FMAP_23_79);
			MULT_80(22)<=signed(DIN_80_7)*signed(FMAP_23_80);
			MULT_81(22)<=signed(DIN_81_7)*signed(FMAP_23_81);
			MULT_82(22)<=signed(DIN_82_7)*signed(FMAP_23_82);
			MULT_83(22)<=signed(DIN_83_7)*signed(FMAP_23_83);
			MULT_84(22)<=signed(DIN_84_7)*signed(FMAP_23_84);
			MULT_85(22)<=signed(DIN_85_7)*signed(FMAP_23_85);
			MULT_86(22)<=signed(DIN_86_7)*signed(FMAP_23_86);
			MULT_87(22)<=signed(DIN_87_7)*signed(FMAP_23_87);
			MULT_88(22)<=signed(DIN_88_7)*signed(FMAP_23_88);
			MULT_89(22)<=signed(DIN_89_7)*signed(FMAP_23_89);
			MULT_90(22)<=signed(DIN_90_7)*signed(FMAP_23_90);
			MULT_91(22)<=signed(DIN_91_7)*signed(FMAP_23_91);
			MULT_92(22)<=signed(DIN_92_7)*signed(FMAP_23_92);
			MULT_93(22)<=signed(DIN_93_7)*signed(FMAP_23_93);
			MULT_94(22)<=signed(DIN_94_7)*signed(FMAP_23_94);
			MULT_95(22)<=signed(DIN_95_7)*signed(FMAP_23_95);
			MULT_96(22)<=signed(DIN_96_7)*signed(FMAP_23_96);
			MULT_97(22)<=signed(DIN_97_7)*signed(FMAP_23_97);
			MULT_98(22)<=signed(DIN_98_7)*signed(FMAP_23_98);
			MULT_99(22)<=signed(DIN_99_7)*signed(FMAP_23_99);
			MULT_100(22)<=signed(DIN_100_7)*signed(FMAP_23_100);
			MULT_101(22)<=signed(DIN_101_7)*signed(FMAP_23_101);
			MULT_102(22)<=signed(DIN_102_7)*signed(FMAP_23_102);
			MULT_103(22)<=signed(DIN_103_7)*signed(FMAP_23_103);
			MULT_104(22)<=signed(DIN_104_7)*signed(FMAP_23_104);
			MULT_105(22)<=signed(DIN_105_7)*signed(FMAP_23_105);
			MULT_106(22)<=signed(DIN_106_7)*signed(FMAP_23_106);
			MULT_107(22)<=signed(DIN_107_7)*signed(FMAP_23_107);
			MULT_108(22)<=signed(DIN_108_7)*signed(FMAP_23_108);
			MULT_109(22)<=signed(DIN_109_7)*signed(FMAP_23_109);
			MULT_110(22)<=signed(DIN_110_7)*signed(FMAP_23_110);
			MULT_111(22)<=signed(DIN_111_7)*signed(FMAP_23_111);
			MULT_112(22)<=signed(DIN_112_7)*signed(FMAP_23_112);
			MULT_113(22)<=signed(DIN_113_7)*signed(FMAP_23_113);
			MULT_114(22)<=signed(DIN_114_7)*signed(FMAP_23_114);
			MULT_115(22)<=signed(DIN_115_7)*signed(FMAP_23_115);
			MULT_116(22)<=signed(DIN_116_7)*signed(FMAP_23_116);
			MULT_117(22)<=signed(DIN_117_7)*signed(FMAP_23_117);
			MULT_118(22)<=signed(DIN_118_7)*signed(FMAP_23_118);
			MULT_119(22)<=signed(DIN_119_7)*signed(FMAP_23_119);
			MULT_120(22)<=signed(DIN_120_7)*signed(FMAP_23_120);

			MULT_1(23)<=signed(DIN_1_7)*signed(FMAP_24_1);
			MULT_2(23)<=signed(DIN_2_7)*signed(FMAP_24_2);
			MULT_3(23)<=signed(DIN_3_7)*signed(FMAP_24_3);
			MULT_4(23)<=signed(DIN_4_7)*signed(FMAP_24_4);
			MULT_5(23)<=signed(DIN_5_7)*signed(FMAP_24_5);
			MULT_6(23)<=signed(DIN_6_7)*signed(FMAP_24_6);
			MULT_7(23)<=signed(DIN_7_7)*signed(FMAP_24_7);
			MULT_8(23)<=signed(DIN_8_7)*signed(FMAP_24_8);
			MULT_9(23)<=signed(DIN_9_7)*signed(FMAP_24_9);
			MULT_10(23)<=signed(DIN_10_7)*signed(FMAP_24_10);
			MULT_11(23)<=signed(DIN_11_7)*signed(FMAP_24_11);
			MULT_12(23)<=signed(DIN_12_7)*signed(FMAP_24_12);
			MULT_13(23)<=signed(DIN_13_7)*signed(FMAP_24_13);
			MULT_14(23)<=signed(DIN_14_7)*signed(FMAP_24_14);
			MULT_15(23)<=signed(DIN_15_7)*signed(FMAP_24_15);
			MULT_16(23)<=signed(DIN_16_7)*signed(FMAP_24_16);
			MULT_17(23)<=signed(DIN_17_7)*signed(FMAP_24_17);
			MULT_18(23)<=signed(DIN_18_7)*signed(FMAP_24_18);
			MULT_19(23)<=signed(DIN_19_7)*signed(FMAP_24_19);
			MULT_20(23)<=signed(DIN_20_7)*signed(FMAP_24_20);
			MULT_21(23)<=signed(DIN_21_7)*signed(FMAP_24_21);
			MULT_22(23)<=signed(DIN_22_7)*signed(FMAP_24_22);
			MULT_23(23)<=signed(DIN_23_7)*signed(FMAP_24_23);
			MULT_24(23)<=signed(DIN_24_7)*signed(FMAP_24_24);
			MULT_25(23)<=signed(DIN_25_7)*signed(FMAP_24_25);
			MULT_26(23)<=signed(DIN_26_7)*signed(FMAP_24_26);
			MULT_27(23)<=signed(DIN_27_7)*signed(FMAP_24_27);
			MULT_28(23)<=signed(DIN_28_7)*signed(FMAP_24_28);
			MULT_29(23)<=signed(DIN_29_7)*signed(FMAP_24_29);
			MULT_30(23)<=signed(DIN_30_7)*signed(FMAP_24_30);
			MULT_31(23)<=signed(DIN_31_7)*signed(FMAP_24_31);
			MULT_32(23)<=signed(DIN_32_7)*signed(FMAP_24_32);
			MULT_33(23)<=signed(DIN_33_7)*signed(FMAP_24_33);
			MULT_34(23)<=signed(DIN_34_7)*signed(FMAP_24_34);
			MULT_35(23)<=signed(DIN_35_7)*signed(FMAP_24_35);
			MULT_36(23)<=signed(DIN_36_7)*signed(FMAP_24_36);
			MULT_37(23)<=signed(DIN_37_7)*signed(FMAP_24_37);
			MULT_38(23)<=signed(DIN_38_7)*signed(FMAP_24_38);
			MULT_39(23)<=signed(DIN_39_7)*signed(FMAP_24_39);
			MULT_40(23)<=signed(DIN_40_7)*signed(FMAP_24_40);
			MULT_41(23)<=signed(DIN_41_7)*signed(FMAP_24_41);
			MULT_42(23)<=signed(DIN_42_7)*signed(FMAP_24_42);
			MULT_43(23)<=signed(DIN_43_7)*signed(FMAP_24_43);
			MULT_44(23)<=signed(DIN_44_7)*signed(FMAP_24_44);
			MULT_45(23)<=signed(DIN_45_7)*signed(FMAP_24_45);
			MULT_46(23)<=signed(DIN_46_7)*signed(FMAP_24_46);
			MULT_47(23)<=signed(DIN_47_7)*signed(FMAP_24_47);
			MULT_48(23)<=signed(DIN_48_7)*signed(FMAP_24_48);
			MULT_49(23)<=signed(DIN_49_7)*signed(FMAP_24_49);
			MULT_50(23)<=signed(DIN_50_7)*signed(FMAP_24_50);
			MULT_51(23)<=signed(DIN_51_7)*signed(FMAP_24_51);
			MULT_52(23)<=signed(DIN_52_7)*signed(FMAP_24_52);
			MULT_53(23)<=signed(DIN_53_7)*signed(FMAP_24_53);
			MULT_54(23)<=signed(DIN_54_7)*signed(FMAP_24_54);
			MULT_55(23)<=signed(DIN_55_7)*signed(FMAP_24_55);
			MULT_56(23)<=signed(DIN_56_7)*signed(FMAP_24_56);
			MULT_57(23)<=signed(DIN_57_7)*signed(FMAP_24_57);
			MULT_58(23)<=signed(DIN_58_7)*signed(FMAP_24_58);
			MULT_59(23)<=signed(DIN_59_7)*signed(FMAP_24_59);
			MULT_60(23)<=signed(DIN_60_7)*signed(FMAP_24_60);
			MULT_61(23)<=signed(DIN_61_7)*signed(FMAP_24_61);
			MULT_62(23)<=signed(DIN_62_7)*signed(FMAP_24_62);
			MULT_63(23)<=signed(DIN_63_7)*signed(FMAP_24_63);
			MULT_64(23)<=signed(DIN_64_7)*signed(FMAP_24_64);
			MULT_65(23)<=signed(DIN_65_7)*signed(FMAP_24_65);
			MULT_66(23)<=signed(DIN_66_7)*signed(FMAP_24_66);
			MULT_67(23)<=signed(DIN_67_7)*signed(FMAP_24_67);
			MULT_68(23)<=signed(DIN_68_7)*signed(FMAP_24_68);
			MULT_69(23)<=signed(DIN_69_7)*signed(FMAP_24_69);
			MULT_70(23)<=signed(DIN_70_7)*signed(FMAP_24_70);
			MULT_71(23)<=signed(DIN_71_7)*signed(FMAP_24_71);
			MULT_72(23)<=signed(DIN_72_7)*signed(FMAP_24_72);
			MULT_73(23)<=signed(DIN_73_7)*signed(FMAP_24_73);
			MULT_74(23)<=signed(DIN_74_7)*signed(FMAP_24_74);
			MULT_75(23)<=signed(DIN_75_7)*signed(FMAP_24_75);
			MULT_76(23)<=signed(DIN_76_7)*signed(FMAP_24_76);
			MULT_77(23)<=signed(DIN_77_7)*signed(FMAP_24_77);
			MULT_78(23)<=signed(DIN_78_7)*signed(FMAP_24_78);
			MULT_79(23)<=signed(DIN_79_7)*signed(FMAP_24_79);
			MULT_80(23)<=signed(DIN_80_7)*signed(FMAP_24_80);
			MULT_81(23)<=signed(DIN_81_7)*signed(FMAP_24_81);
			MULT_82(23)<=signed(DIN_82_7)*signed(FMAP_24_82);
			MULT_83(23)<=signed(DIN_83_7)*signed(FMAP_24_83);
			MULT_84(23)<=signed(DIN_84_7)*signed(FMAP_24_84);
			MULT_85(23)<=signed(DIN_85_7)*signed(FMAP_24_85);
			MULT_86(23)<=signed(DIN_86_7)*signed(FMAP_24_86);
			MULT_87(23)<=signed(DIN_87_7)*signed(FMAP_24_87);
			MULT_88(23)<=signed(DIN_88_7)*signed(FMAP_24_88);
			MULT_89(23)<=signed(DIN_89_7)*signed(FMAP_24_89);
			MULT_90(23)<=signed(DIN_90_7)*signed(FMAP_24_90);
			MULT_91(23)<=signed(DIN_91_7)*signed(FMAP_24_91);
			MULT_92(23)<=signed(DIN_92_7)*signed(FMAP_24_92);
			MULT_93(23)<=signed(DIN_93_7)*signed(FMAP_24_93);
			MULT_94(23)<=signed(DIN_94_7)*signed(FMAP_24_94);
			MULT_95(23)<=signed(DIN_95_7)*signed(FMAP_24_95);
			MULT_96(23)<=signed(DIN_96_7)*signed(FMAP_24_96);
			MULT_97(23)<=signed(DIN_97_7)*signed(FMAP_24_97);
			MULT_98(23)<=signed(DIN_98_7)*signed(FMAP_24_98);
			MULT_99(23)<=signed(DIN_99_7)*signed(FMAP_24_99);
			MULT_100(23)<=signed(DIN_100_7)*signed(FMAP_24_100);
			MULT_101(23)<=signed(DIN_101_7)*signed(FMAP_24_101);
			MULT_102(23)<=signed(DIN_102_7)*signed(FMAP_24_102);
			MULT_103(23)<=signed(DIN_103_7)*signed(FMAP_24_103);
			MULT_104(23)<=signed(DIN_104_7)*signed(FMAP_24_104);
			MULT_105(23)<=signed(DIN_105_7)*signed(FMAP_24_105);
			MULT_106(23)<=signed(DIN_106_7)*signed(FMAP_24_106);
			MULT_107(23)<=signed(DIN_107_7)*signed(FMAP_24_107);
			MULT_108(23)<=signed(DIN_108_7)*signed(FMAP_24_108);
			MULT_109(23)<=signed(DIN_109_7)*signed(FMAP_24_109);
			MULT_110(23)<=signed(DIN_110_7)*signed(FMAP_24_110);
			MULT_111(23)<=signed(DIN_111_7)*signed(FMAP_24_111);
			MULT_112(23)<=signed(DIN_112_7)*signed(FMAP_24_112);
			MULT_113(23)<=signed(DIN_113_7)*signed(FMAP_24_113);
			MULT_114(23)<=signed(DIN_114_7)*signed(FMAP_24_114);
			MULT_115(23)<=signed(DIN_115_7)*signed(FMAP_24_115);
			MULT_116(23)<=signed(DIN_116_7)*signed(FMAP_24_116);
			MULT_117(23)<=signed(DIN_117_7)*signed(FMAP_24_117);
			MULT_118(23)<=signed(DIN_118_7)*signed(FMAP_24_118);
			MULT_119(23)<=signed(DIN_119_7)*signed(FMAP_24_119);
			MULT_120(23)<=signed(DIN_120_7)*signed(FMAP_24_120);

			MULT_1(24)<=signed(DIN_1_7)*signed(FMAP_25_1);
			MULT_2(24)<=signed(DIN_2_7)*signed(FMAP_25_2);
			MULT_3(24)<=signed(DIN_3_7)*signed(FMAP_25_3);
			MULT_4(24)<=signed(DIN_4_7)*signed(FMAP_25_4);
			MULT_5(24)<=signed(DIN_5_7)*signed(FMAP_25_5);
			MULT_6(24)<=signed(DIN_6_7)*signed(FMAP_25_6);
			MULT_7(24)<=signed(DIN_7_7)*signed(FMAP_25_7);
			MULT_8(24)<=signed(DIN_8_7)*signed(FMAP_25_8);
			MULT_9(24)<=signed(DIN_9_7)*signed(FMAP_25_9);
			MULT_10(24)<=signed(DIN_10_7)*signed(FMAP_25_10);
			MULT_11(24)<=signed(DIN_11_7)*signed(FMAP_25_11);
			MULT_12(24)<=signed(DIN_12_7)*signed(FMAP_25_12);
			MULT_13(24)<=signed(DIN_13_7)*signed(FMAP_25_13);
			MULT_14(24)<=signed(DIN_14_7)*signed(FMAP_25_14);
			MULT_15(24)<=signed(DIN_15_7)*signed(FMAP_25_15);
			MULT_16(24)<=signed(DIN_16_7)*signed(FMAP_25_16);
			MULT_17(24)<=signed(DIN_17_7)*signed(FMAP_25_17);
			MULT_18(24)<=signed(DIN_18_7)*signed(FMAP_25_18);
			MULT_19(24)<=signed(DIN_19_7)*signed(FMAP_25_19);
			MULT_20(24)<=signed(DIN_20_7)*signed(FMAP_25_20);
			MULT_21(24)<=signed(DIN_21_7)*signed(FMAP_25_21);
			MULT_22(24)<=signed(DIN_22_7)*signed(FMAP_25_22);
			MULT_23(24)<=signed(DIN_23_7)*signed(FMAP_25_23);
			MULT_24(24)<=signed(DIN_24_7)*signed(FMAP_25_24);
			MULT_25(24)<=signed(DIN_25_7)*signed(FMAP_25_25);
			MULT_26(24)<=signed(DIN_26_7)*signed(FMAP_25_26);
			MULT_27(24)<=signed(DIN_27_7)*signed(FMAP_25_27);
			MULT_28(24)<=signed(DIN_28_7)*signed(FMAP_25_28);
			MULT_29(24)<=signed(DIN_29_7)*signed(FMAP_25_29);
			MULT_30(24)<=signed(DIN_30_7)*signed(FMAP_25_30);
			MULT_31(24)<=signed(DIN_31_7)*signed(FMAP_25_31);
			MULT_32(24)<=signed(DIN_32_7)*signed(FMAP_25_32);
			MULT_33(24)<=signed(DIN_33_7)*signed(FMAP_25_33);
			MULT_34(24)<=signed(DIN_34_7)*signed(FMAP_25_34);
			MULT_35(24)<=signed(DIN_35_7)*signed(FMAP_25_35);
			MULT_36(24)<=signed(DIN_36_7)*signed(FMAP_25_36);
			MULT_37(24)<=signed(DIN_37_7)*signed(FMAP_25_37);
			MULT_38(24)<=signed(DIN_38_7)*signed(FMAP_25_38);
			MULT_39(24)<=signed(DIN_39_7)*signed(FMAP_25_39);
			MULT_40(24)<=signed(DIN_40_7)*signed(FMAP_25_40);
			MULT_41(24)<=signed(DIN_41_7)*signed(FMAP_25_41);
			MULT_42(24)<=signed(DIN_42_7)*signed(FMAP_25_42);
			MULT_43(24)<=signed(DIN_43_7)*signed(FMAP_25_43);
			MULT_44(24)<=signed(DIN_44_7)*signed(FMAP_25_44);
			MULT_45(24)<=signed(DIN_45_7)*signed(FMAP_25_45);
			MULT_46(24)<=signed(DIN_46_7)*signed(FMAP_25_46);
			MULT_47(24)<=signed(DIN_47_7)*signed(FMAP_25_47);
			MULT_48(24)<=signed(DIN_48_7)*signed(FMAP_25_48);
			MULT_49(24)<=signed(DIN_49_7)*signed(FMAP_25_49);
			MULT_50(24)<=signed(DIN_50_7)*signed(FMAP_25_50);
			MULT_51(24)<=signed(DIN_51_7)*signed(FMAP_25_51);
			MULT_52(24)<=signed(DIN_52_7)*signed(FMAP_25_52);
			MULT_53(24)<=signed(DIN_53_7)*signed(FMAP_25_53);
			MULT_54(24)<=signed(DIN_54_7)*signed(FMAP_25_54);
			MULT_55(24)<=signed(DIN_55_7)*signed(FMAP_25_55);
			MULT_56(24)<=signed(DIN_56_7)*signed(FMAP_25_56);
			MULT_57(24)<=signed(DIN_57_7)*signed(FMAP_25_57);
			MULT_58(24)<=signed(DIN_58_7)*signed(FMAP_25_58);
			MULT_59(24)<=signed(DIN_59_7)*signed(FMAP_25_59);
			MULT_60(24)<=signed(DIN_60_7)*signed(FMAP_25_60);
			MULT_61(24)<=signed(DIN_61_7)*signed(FMAP_25_61);
			MULT_62(24)<=signed(DIN_62_7)*signed(FMAP_25_62);
			MULT_63(24)<=signed(DIN_63_7)*signed(FMAP_25_63);
			MULT_64(24)<=signed(DIN_64_7)*signed(FMAP_25_64);
			MULT_65(24)<=signed(DIN_65_7)*signed(FMAP_25_65);
			MULT_66(24)<=signed(DIN_66_7)*signed(FMAP_25_66);
			MULT_67(24)<=signed(DIN_67_7)*signed(FMAP_25_67);
			MULT_68(24)<=signed(DIN_68_7)*signed(FMAP_25_68);
			MULT_69(24)<=signed(DIN_69_7)*signed(FMAP_25_69);
			MULT_70(24)<=signed(DIN_70_7)*signed(FMAP_25_70);
			MULT_71(24)<=signed(DIN_71_7)*signed(FMAP_25_71);
			MULT_72(24)<=signed(DIN_72_7)*signed(FMAP_25_72);
			MULT_73(24)<=signed(DIN_73_7)*signed(FMAP_25_73);
			MULT_74(24)<=signed(DIN_74_7)*signed(FMAP_25_74);
			MULT_75(24)<=signed(DIN_75_7)*signed(FMAP_25_75);
			MULT_76(24)<=signed(DIN_76_7)*signed(FMAP_25_76);
			MULT_77(24)<=signed(DIN_77_7)*signed(FMAP_25_77);
			MULT_78(24)<=signed(DIN_78_7)*signed(FMAP_25_78);
			MULT_79(24)<=signed(DIN_79_7)*signed(FMAP_25_79);
			MULT_80(24)<=signed(DIN_80_7)*signed(FMAP_25_80);
			MULT_81(24)<=signed(DIN_81_7)*signed(FMAP_25_81);
			MULT_82(24)<=signed(DIN_82_7)*signed(FMAP_25_82);
			MULT_83(24)<=signed(DIN_83_7)*signed(FMAP_25_83);
			MULT_84(24)<=signed(DIN_84_7)*signed(FMAP_25_84);
			MULT_85(24)<=signed(DIN_85_7)*signed(FMAP_25_85);
			MULT_86(24)<=signed(DIN_86_7)*signed(FMAP_25_86);
			MULT_87(24)<=signed(DIN_87_7)*signed(FMAP_25_87);
			MULT_88(24)<=signed(DIN_88_7)*signed(FMAP_25_88);
			MULT_89(24)<=signed(DIN_89_7)*signed(FMAP_25_89);
			MULT_90(24)<=signed(DIN_90_7)*signed(FMAP_25_90);
			MULT_91(24)<=signed(DIN_91_7)*signed(FMAP_25_91);
			MULT_92(24)<=signed(DIN_92_7)*signed(FMAP_25_92);
			MULT_93(24)<=signed(DIN_93_7)*signed(FMAP_25_93);
			MULT_94(24)<=signed(DIN_94_7)*signed(FMAP_25_94);
			MULT_95(24)<=signed(DIN_95_7)*signed(FMAP_25_95);
			MULT_96(24)<=signed(DIN_96_7)*signed(FMAP_25_96);
			MULT_97(24)<=signed(DIN_97_7)*signed(FMAP_25_97);
			MULT_98(24)<=signed(DIN_98_7)*signed(FMAP_25_98);
			MULT_99(24)<=signed(DIN_99_7)*signed(FMAP_25_99);
			MULT_100(24)<=signed(DIN_100_7)*signed(FMAP_25_100);
			MULT_101(24)<=signed(DIN_101_7)*signed(FMAP_25_101);
			MULT_102(24)<=signed(DIN_102_7)*signed(FMAP_25_102);
			MULT_103(24)<=signed(DIN_103_7)*signed(FMAP_25_103);
			MULT_104(24)<=signed(DIN_104_7)*signed(FMAP_25_104);
			MULT_105(24)<=signed(DIN_105_7)*signed(FMAP_25_105);
			MULT_106(24)<=signed(DIN_106_7)*signed(FMAP_25_106);
			MULT_107(24)<=signed(DIN_107_7)*signed(FMAP_25_107);
			MULT_108(24)<=signed(DIN_108_7)*signed(FMAP_25_108);
			MULT_109(24)<=signed(DIN_109_7)*signed(FMAP_25_109);
			MULT_110(24)<=signed(DIN_110_7)*signed(FMAP_25_110);
			MULT_111(24)<=signed(DIN_111_7)*signed(FMAP_25_111);
			MULT_112(24)<=signed(DIN_112_7)*signed(FMAP_25_112);
			MULT_113(24)<=signed(DIN_113_7)*signed(FMAP_25_113);
			MULT_114(24)<=signed(DIN_114_7)*signed(FMAP_25_114);
			MULT_115(24)<=signed(DIN_115_7)*signed(FMAP_25_115);
			MULT_116(24)<=signed(DIN_116_7)*signed(FMAP_25_116);
			MULT_117(24)<=signed(DIN_117_7)*signed(FMAP_25_117);
			MULT_118(24)<=signed(DIN_118_7)*signed(FMAP_25_118);
			MULT_119(24)<=signed(DIN_119_7)*signed(FMAP_25_119);
			MULT_120(24)<=signed(DIN_120_7)*signed(FMAP_25_120);

			MULT_1(25)<=signed(DIN_1_7)*signed(FMAP_26_1);
			MULT_2(25)<=signed(DIN_2_7)*signed(FMAP_26_2);
			MULT_3(25)<=signed(DIN_3_7)*signed(FMAP_26_3);
			MULT_4(25)<=signed(DIN_4_7)*signed(FMAP_26_4);
			MULT_5(25)<=signed(DIN_5_7)*signed(FMAP_26_5);
			MULT_6(25)<=signed(DIN_6_7)*signed(FMAP_26_6);
			MULT_7(25)<=signed(DIN_7_7)*signed(FMAP_26_7);
			MULT_8(25)<=signed(DIN_8_7)*signed(FMAP_26_8);
			MULT_9(25)<=signed(DIN_9_7)*signed(FMAP_26_9);
			MULT_10(25)<=signed(DIN_10_7)*signed(FMAP_26_10);
			MULT_11(25)<=signed(DIN_11_7)*signed(FMAP_26_11);
			MULT_12(25)<=signed(DIN_12_7)*signed(FMAP_26_12);
			MULT_13(25)<=signed(DIN_13_7)*signed(FMAP_26_13);
			MULT_14(25)<=signed(DIN_14_7)*signed(FMAP_26_14);
			MULT_15(25)<=signed(DIN_15_7)*signed(FMAP_26_15);
			MULT_16(25)<=signed(DIN_16_7)*signed(FMAP_26_16);
			MULT_17(25)<=signed(DIN_17_7)*signed(FMAP_26_17);
			MULT_18(25)<=signed(DIN_18_7)*signed(FMAP_26_18);
			MULT_19(25)<=signed(DIN_19_7)*signed(FMAP_26_19);
			MULT_20(25)<=signed(DIN_20_7)*signed(FMAP_26_20);
			MULT_21(25)<=signed(DIN_21_7)*signed(FMAP_26_21);
			MULT_22(25)<=signed(DIN_22_7)*signed(FMAP_26_22);
			MULT_23(25)<=signed(DIN_23_7)*signed(FMAP_26_23);
			MULT_24(25)<=signed(DIN_24_7)*signed(FMAP_26_24);
			MULT_25(25)<=signed(DIN_25_7)*signed(FMAP_26_25);
			MULT_26(25)<=signed(DIN_26_7)*signed(FMAP_26_26);
			MULT_27(25)<=signed(DIN_27_7)*signed(FMAP_26_27);
			MULT_28(25)<=signed(DIN_28_7)*signed(FMAP_26_28);
			MULT_29(25)<=signed(DIN_29_7)*signed(FMAP_26_29);
			MULT_30(25)<=signed(DIN_30_7)*signed(FMAP_26_30);
			MULT_31(25)<=signed(DIN_31_7)*signed(FMAP_26_31);
			MULT_32(25)<=signed(DIN_32_7)*signed(FMAP_26_32);
			MULT_33(25)<=signed(DIN_33_7)*signed(FMAP_26_33);
			MULT_34(25)<=signed(DIN_34_7)*signed(FMAP_26_34);
			MULT_35(25)<=signed(DIN_35_7)*signed(FMAP_26_35);
			MULT_36(25)<=signed(DIN_36_7)*signed(FMAP_26_36);
			MULT_37(25)<=signed(DIN_37_7)*signed(FMAP_26_37);
			MULT_38(25)<=signed(DIN_38_7)*signed(FMAP_26_38);
			MULT_39(25)<=signed(DIN_39_7)*signed(FMAP_26_39);
			MULT_40(25)<=signed(DIN_40_7)*signed(FMAP_26_40);
			MULT_41(25)<=signed(DIN_41_7)*signed(FMAP_26_41);
			MULT_42(25)<=signed(DIN_42_7)*signed(FMAP_26_42);
			MULT_43(25)<=signed(DIN_43_7)*signed(FMAP_26_43);
			MULT_44(25)<=signed(DIN_44_7)*signed(FMAP_26_44);
			MULT_45(25)<=signed(DIN_45_7)*signed(FMAP_26_45);
			MULT_46(25)<=signed(DIN_46_7)*signed(FMAP_26_46);
			MULT_47(25)<=signed(DIN_47_7)*signed(FMAP_26_47);
			MULT_48(25)<=signed(DIN_48_7)*signed(FMAP_26_48);
			MULT_49(25)<=signed(DIN_49_7)*signed(FMAP_26_49);
			MULT_50(25)<=signed(DIN_50_7)*signed(FMAP_26_50);
			MULT_51(25)<=signed(DIN_51_7)*signed(FMAP_26_51);
			MULT_52(25)<=signed(DIN_52_7)*signed(FMAP_26_52);
			MULT_53(25)<=signed(DIN_53_7)*signed(FMAP_26_53);
			MULT_54(25)<=signed(DIN_54_7)*signed(FMAP_26_54);
			MULT_55(25)<=signed(DIN_55_7)*signed(FMAP_26_55);
			MULT_56(25)<=signed(DIN_56_7)*signed(FMAP_26_56);
			MULT_57(25)<=signed(DIN_57_7)*signed(FMAP_26_57);
			MULT_58(25)<=signed(DIN_58_7)*signed(FMAP_26_58);
			MULT_59(25)<=signed(DIN_59_7)*signed(FMAP_26_59);
			MULT_60(25)<=signed(DIN_60_7)*signed(FMAP_26_60);
			MULT_61(25)<=signed(DIN_61_7)*signed(FMAP_26_61);
			MULT_62(25)<=signed(DIN_62_7)*signed(FMAP_26_62);
			MULT_63(25)<=signed(DIN_63_7)*signed(FMAP_26_63);
			MULT_64(25)<=signed(DIN_64_7)*signed(FMAP_26_64);
			MULT_65(25)<=signed(DIN_65_7)*signed(FMAP_26_65);
			MULT_66(25)<=signed(DIN_66_7)*signed(FMAP_26_66);
			MULT_67(25)<=signed(DIN_67_7)*signed(FMAP_26_67);
			MULT_68(25)<=signed(DIN_68_7)*signed(FMAP_26_68);
			MULT_69(25)<=signed(DIN_69_7)*signed(FMAP_26_69);
			MULT_70(25)<=signed(DIN_70_7)*signed(FMAP_26_70);
			MULT_71(25)<=signed(DIN_71_7)*signed(FMAP_26_71);
			MULT_72(25)<=signed(DIN_72_7)*signed(FMAP_26_72);
			MULT_73(25)<=signed(DIN_73_7)*signed(FMAP_26_73);
			MULT_74(25)<=signed(DIN_74_7)*signed(FMAP_26_74);
			MULT_75(25)<=signed(DIN_75_7)*signed(FMAP_26_75);
			MULT_76(25)<=signed(DIN_76_7)*signed(FMAP_26_76);
			MULT_77(25)<=signed(DIN_77_7)*signed(FMAP_26_77);
			MULT_78(25)<=signed(DIN_78_7)*signed(FMAP_26_78);
			MULT_79(25)<=signed(DIN_79_7)*signed(FMAP_26_79);
			MULT_80(25)<=signed(DIN_80_7)*signed(FMAP_26_80);
			MULT_81(25)<=signed(DIN_81_7)*signed(FMAP_26_81);
			MULT_82(25)<=signed(DIN_82_7)*signed(FMAP_26_82);
			MULT_83(25)<=signed(DIN_83_7)*signed(FMAP_26_83);
			MULT_84(25)<=signed(DIN_84_7)*signed(FMAP_26_84);
			MULT_85(25)<=signed(DIN_85_7)*signed(FMAP_26_85);
			MULT_86(25)<=signed(DIN_86_7)*signed(FMAP_26_86);
			MULT_87(25)<=signed(DIN_87_7)*signed(FMAP_26_87);
			MULT_88(25)<=signed(DIN_88_7)*signed(FMAP_26_88);
			MULT_89(25)<=signed(DIN_89_7)*signed(FMAP_26_89);
			MULT_90(25)<=signed(DIN_90_7)*signed(FMAP_26_90);
			MULT_91(25)<=signed(DIN_91_7)*signed(FMAP_26_91);
			MULT_92(25)<=signed(DIN_92_7)*signed(FMAP_26_92);
			MULT_93(25)<=signed(DIN_93_7)*signed(FMAP_26_93);
			MULT_94(25)<=signed(DIN_94_7)*signed(FMAP_26_94);
			MULT_95(25)<=signed(DIN_95_7)*signed(FMAP_26_95);
			MULT_96(25)<=signed(DIN_96_7)*signed(FMAP_26_96);
			MULT_97(25)<=signed(DIN_97_7)*signed(FMAP_26_97);
			MULT_98(25)<=signed(DIN_98_7)*signed(FMAP_26_98);
			MULT_99(25)<=signed(DIN_99_7)*signed(FMAP_26_99);
			MULT_100(25)<=signed(DIN_100_7)*signed(FMAP_26_100);
			MULT_101(25)<=signed(DIN_101_7)*signed(FMAP_26_101);
			MULT_102(25)<=signed(DIN_102_7)*signed(FMAP_26_102);
			MULT_103(25)<=signed(DIN_103_7)*signed(FMAP_26_103);
			MULT_104(25)<=signed(DIN_104_7)*signed(FMAP_26_104);
			MULT_105(25)<=signed(DIN_105_7)*signed(FMAP_26_105);
			MULT_106(25)<=signed(DIN_106_7)*signed(FMAP_26_106);
			MULT_107(25)<=signed(DIN_107_7)*signed(FMAP_26_107);
			MULT_108(25)<=signed(DIN_108_7)*signed(FMAP_26_108);
			MULT_109(25)<=signed(DIN_109_7)*signed(FMAP_26_109);
			MULT_110(25)<=signed(DIN_110_7)*signed(FMAP_26_110);
			MULT_111(25)<=signed(DIN_111_7)*signed(FMAP_26_111);
			MULT_112(25)<=signed(DIN_112_7)*signed(FMAP_26_112);
			MULT_113(25)<=signed(DIN_113_7)*signed(FMAP_26_113);
			MULT_114(25)<=signed(DIN_114_7)*signed(FMAP_26_114);
			MULT_115(25)<=signed(DIN_115_7)*signed(FMAP_26_115);
			MULT_116(25)<=signed(DIN_116_7)*signed(FMAP_26_116);
			MULT_117(25)<=signed(DIN_117_7)*signed(FMAP_26_117);
			MULT_118(25)<=signed(DIN_118_7)*signed(FMAP_26_118);
			MULT_119(25)<=signed(DIN_119_7)*signed(FMAP_26_119);
			MULT_120(25)<=signed(DIN_120_7)*signed(FMAP_26_120);

			MULT_1(26)<=signed(DIN_1_7)*signed(FMAP_27_1);
			MULT_2(26)<=signed(DIN_2_7)*signed(FMAP_27_2);
			MULT_3(26)<=signed(DIN_3_7)*signed(FMAP_27_3);
			MULT_4(26)<=signed(DIN_4_7)*signed(FMAP_27_4);
			MULT_5(26)<=signed(DIN_5_7)*signed(FMAP_27_5);
			MULT_6(26)<=signed(DIN_6_7)*signed(FMAP_27_6);
			MULT_7(26)<=signed(DIN_7_7)*signed(FMAP_27_7);
			MULT_8(26)<=signed(DIN_8_7)*signed(FMAP_27_8);
			MULT_9(26)<=signed(DIN_9_7)*signed(FMAP_27_9);
			MULT_10(26)<=signed(DIN_10_7)*signed(FMAP_27_10);
			MULT_11(26)<=signed(DIN_11_7)*signed(FMAP_27_11);
			MULT_12(26)<=signed(DIN_12_7)*signed(FMAP_27_12);
			MULT_13(26)<=signed(DIN_13_7)*signed(FMAP_27_13);
			MULT_14(26)<=signed(DIN_14_7)*signed(FMAP_27_14);
			MULT_15(26)<=signed(DIN_15_7)*signed(FMAP_27_15);
			MULT_16(26)<=signed(DIN_16_7)*signed(FMAP_27_16);
			MULT_17(26)<=signed(DIN_17_7)*signed(FMAP_27_17);
			MULT_18(26)<=signed(DIN_18_7)*signed(FMAP_27_18);
			MULT_19(26)<=signed(DIN_19_7)*signed(FMAP_27_19);
			MULT_20(26)<=signed(DIN_20_7)*signed(FMAP_27_20);
			MULT_21(26)<=signed(DIN_21_7)*signed(FMAP_27_21);
			MULT_22(26)<=signed(DIN_22_7)*signed(FMAP_27_22);
			MULT_23(26)<=signed(DIN_23_7)*signed(FMAP_27_23);
			MULT_24(26)<=signed(DIN_24_7)*signed(FMAP_27_24);
			MULT_25(26)<=signed(DIN_25_7)*signed(FMAP_27_25);
			MULT_26(26)<=signed(DIN_26_7)*signed(FMAP_27_26);
			MULT_27(26)<=signed(DIN_27_7)*signed(FMAP_27_27);
			MULT_28(26)<=signed(DIN_28_7)*signed(FMAP_27_28);
			MULT_29(26)<=signed(DIN_29_7)*signed(FMAP_27_29);
			MULT_30(26)<=signed(DIN_30_7)*signed(FMAP_27_30);
			MULT_31(26)<=signed(DIN_31_7)*signed(FMAP_27_31);
			MULT_32(26)<=signed(DIN_32_7)*signed(FMAP_27_32);
			MULT_33(26)<=signed(DIN_33_7)*signed(FMAP_27_33);
			MULT_34(26)<=signed(DIN_34_7)*signed(FMAP_27_34);
			MULT_35(26)<=signed(DIN_35_7)*signed(FMAP_27_35);
			MULT_36(26)<=signed(DIN_36_7)*signed(FMAP_27_36);
			MULT_37(26)<=signed(DIN_37_7)*signed(FMAP_27_37);
			MULT_38(26)<=signed(DIN_38_7)*signed(FMAP_27_38);
			MULT_39(26)<=signed(DIN_39_7)*signed(FMAP_27_39);
			MULT_40(26)<=signed(DIN_40_7)*signed(FMAP_27_40);
			MULT_41(26)<=signed(DIN_41_7)*signed(FMAP_27_41);
			MULT_42(26)<=signed(DIN_42_7)*signed(FMAP_27_42);
			MULT_43(26)<=signed(DIN_43_7)*signed(FMAP_27_43);
			MULT_44(26)<=signed(DIN_44_7)*signed(FMAP_27_44);
			MULT_45(26)<=signed(DIN_45_7)*signed(FMAP_27_45);
			MULT_46(26)<=signed(DIN_46_7)*signed(FMAP_27_46);
			MULT_47(26)<=signed(DIN_47_7)*signed(FMAP_27_47);
			MULT_48(26)<=signed(DIN_48_7)*signed(FMAP_27_48);
			MULT_49(26)<=signed(DIN_49_7)*signed(FMAP_27_49);
			MULT_50(26)<=signed(DIN_50_7)*signed(FMAP_27_50);
			MULT_51(26)<=signed(DIN_51_7)*signed(FMAP_27_51);
			MULT_52(26)<=signed(DIN_52_7)*signed(FMAP_27_52);
			MULT_53(26)<=signed(DIN_53_7)*signed(FMAP_27_53);
			MULT_54(26)<=signed(DIN_54_7)*signed(FMAP_27_54);
			MULT_55(26)<=signed(DIN_55_7)*signed(FMAP_27_55);
			MULT_56(26)<=signed(DIN_56_7)*signed(FMAP_27_56);
			MULT_57(26)<=signed(DIN_57_7)*signed(FMAP_27_57);
			MULT_58(26)<=signed(DIN_58_7)*signed(FMAP_27_58);
			MULT_59(26)<=signed(DIN_59_7)*signed(FMAP_27_59);
			MULT_60(26)<=signed(DIN_60_7)*signed(FMAP_27_60);
			MULT_61(26)<=signed(DIN_61_7)*signed(FMAP_27_61);
			MULT_62(26)<=signed(DIN_62_7)*signed(FMAP_27_62);
			MULT_63(26)<=signed(DIN_63_7)*signed(FMAP_27_63);
			MULT_64(26)<=signed(DIN_64_7)*signed(FMAP_27_64);
			MULT_65(26)<=signed(DIN_65_7)*signed(FMAP_27_65);
			MULT_66(26)<=signed(DIN_66_7)*signed(FMAP_27_66);
			MULT_67(26)<=signed(DIN_67_7)*signed(FMAP_27_67);
			MULT_68(26)<=signed(DIN_68_7)*signed(FMAP_27_68);
			MULT_69(26)<=signed(DIN_69_7)*signed(FMAP_27_69);
			MULT_70(26)<=signed(DIN_70_7)*signed(FMAP_27_70);
			MULT_71(26)<=signed(DIN_71_7)*signed(FMAP_27_71);
			MULT_72(26)<=signed(DIN_72_7)*signed(FMAP_27_72);
			MULT_73(26)<=signed(DIN_73_7)*signed(FMAP_27_73);
			MULT_74(26)<=signed(DIN_74_7)*signed(FMAP_27_74);
			MULT_75(26)<=signed(DIN_75_7)*signed(FMAP_27_75);
			MULT_76(26)<=signed(DIN_76_7)*signed(FMAP_27_76);
			MULT_77(26)<=signed(DIN_77_7)*signed(FMAP_27_77);
			MULT_78(26)<=signed(DIN_78_7)*signed(FMAP_27_78);
			MULT_79(26)<=signed(DIN_79_7)*signed(FMAP_27_79);
			MULT_80(26)<=signed(DIN_80_7)*signed(FMAP_27_80);
			MULT_81(26)<=signed(DIN_81_7)*signed(FMAP_27_81);
			MULT_82(26)<=signed(DIN_82_7)*signed(FMAP_27_82);
			MULT_83(26)<=signed(DIN_83_7)*signed(FMAP_27_83);
			MULT_84(26)<=signed(DIN_84_7)*signed(FMAP_27_84);
			MULT_85(26)<=signed(DIN_85_7)*signed(FMAP_27_85);
			MULT_86(26)<=signed(DIN_86_7)*signed(FMAP_27_86);
			MULT_87(26)<=signed(DIN_87_7)*signed(FMAP_27_87);
			MULT_88(26)<=signed(DIN_88_7)*signed(FMAP_27_88);
			MULT_89(26)<=signed(DIN_89_7)*signed(FMAP_27_89);
			MULT_90(26)<=signed(DIN_90_7)*signed(FMAP_27_90);
			MULT_91(26)<=signed(DIN_91_7)*signed(FMAP_27_91);
			MULT_92(26)<=signed(DIN_92_7)*signed(FMAP_27_92);
			MULT_93(26)<=signed(DIN_93_7)*signed(FMAP_27_93);
			MULT_94(26)<=signed(DIN_94_7)*signed(FMAP_27_94);
			MULT_95(26)<=signed(DIN_95_7)*signed(FMAP_27_95);
			MULT_96(26)<=signed(DIN_96_7)*signed(FMAP_27_96);
			MULT_97(26)<=signed(DIN_97_7)*signed(FMAP_27_97);
			MULT_98(26)<=signed(DIN_98_7)*signed(FMAP_27_98);
			MULT_99(26)<=signed(DIN_99_7)*signed(FMAP_27_99);
			MULT_100(26)<=signed(DIN_100_7)*signed(FMAP_27_100);
			MULT_101(26)<=signed(DIN_101_7)*signed(FMAP_27_101);
			MULT_102(26)<=signed(DIN_102_7)*signed(FMAP_27_102);
			MULT_103(26)<=signed(DIN_103_7)*signed(FMAP_27_103);
			MULT_104(26)<=signed(DIN_104_7)*signed(FMAP_27_104);
			MULT_105(26)<=signed(DIN_105_7)*signed(FMAP_27_105);
			MULT_106(26)<=signed(DIN_106_7)*signed(FMAP_27_106);
			MULT_107(26)<=signed(DIN_107_7)*signed(FMAP_27_107);
			MULT_108(26)<=signed(DIN_108_7)*signed(FMAP_27_108);
			MULT_109(26)<=signed(DIN_109_7)*signed(FMAP_27_109);
			MULT_110(26)<=signed(DIN_110_7)*signed(FMAP_27_110);
			MULT_111(26)<=signed(DIN_111_7)*signed(FMAP_27_111);
			MULT_112(26)<=signed(DIN_112_7)*signed(FMAP_27_112);
			MULT_113(26)<=signed(DIN_113_7)*signed(FMAP_27_113);
			MULT_114(26)<=signed(DIN_114_7)*signed(FMAP_27_114);
			MULT_115(26)<=signed(DIN_115_7)*signed(FMAP_27_115);
			MULT_116(26)<=signed(DIN_116_7)*signed(FMAP_27_116);
			MULT_117(26)<=signed(DIN_117_7)*signed(FMAP_27_117);
			MULT_118(26)<=signed(DIN_118_7)*signed(FMAP_27_118);
			MULT_119(26)<=signed(DIN_119_7)*signed(FMAP_27_119);
			MULT_120(26)<=signed(DIN_120_7)*signed(FMAP_27_120);

			MULT_1(27)<=signed(DIN_1_7)*signed(FMAP_28_1);
			MULT_2(27)<=signed(DIN_2_7)*signed(FMAP_28_2);
			MULT_3(27)<=signed(DIN_3_7)*signed(FMAP_28_3);
			MULT_4(27)<=signed(DIN_4_7)*signed(FMAP_28_4);
			MULT_5(27)<=signed(DIN_5_7)*signed(FMAP_28_5);
			MULT_6(27)<=signed(DIN_6_7)*signed(FMAP_28_6);
			MULT_7(27)<=signed(DIN_7_7)*signed(FMAP_28_7);
			MULT_8(27)<=signed(DIN_8_7)*signed(FMAP_28_8);
			MULT_9(27)<=signed(DIN_9_7)*signed(FMAP_28_9);
			MULT_10(27)<=signed(DIN_10_7)*signed(FMAP_28_10);
			MULT_11(27)<=signed(DIN_11_7)*signed(FMAP_28_11);
			MULT_12(27)<=signed(DIN_12_7)*signed(FMAP_28_12);
			MULT_13(27)<=signed(DIN_13_7)*signed(FMAP_28_13);
			MULT_14(27)<=signed(DIN_14_7)*signed(FMAP_28_14);
			MULT_15(27)<=signed(DIN_15_7)*signed(FMAP_28_15);
			MULT_16(27)<=signed(DIN_16_7)*signed(FMAP_28_16);
			MULT_17(27)<=signed(DIN_17_7)*signed(FMAP_28_17);
			MULT_18(27)<=signed(DIN_18_7)*signed(FMAP_28_18);
			MULT_19(27)<=signed(DIN_19_7)*signed(FMAP_28_19);
			MULT_20(27)<=signed(DIN_20_7)*signed(FMAP_28_20);
			MULT_21(27)<=signed(DIN_21_7)*signed(FMAP_28_21);
			MULT_22(27)<=signed(DIN_22_7)*signed(FMAP_28_22);
			MULT_23(27)<=signed(DIN_23_7)*signed(FMAP_28_23);
			MULT_24(27)<=signed(DIN_24_7)*signed(FMAP_28_24);
			MULT_25(27)<=signed(DIN_25_7)*signed(FMAP_28_25);
			MULT_26(27)<=signed(DIN_26_7)*signed(FMAP_28_26);
			MULT_27(27)<=signed(DIN_27_7)*signed(FMAP_28_27);
			MULT_28(27)<=signed(DIN_28_7)*signed(FMAP_28_28);
			MULT_29(27)<=signed(DIN_29_7)*signed(FMAP_28_29);
			MULT_30(27)<=signed(DIN_30_7)*signed(FMAP_28_30);
			MULT_31(27)<=signed(DIN_31_7)*signed(FMAP_28_31);
			MULT_32(27)<=signed(DIN_32_7)*signed(FMAP_28_32);
			MULT_33(27)<=signed(DIN_33_7)*signed(FMAP_28_33);
			MULT_34(27)<=signed(DIN_34_7)*signed(FMAP_28_34);
			MULT_35(27)<=signed(DIN_35_7)*signed(FMAP_28_35);
			MULT_36(27)<=signed(DIN_36_7)*signed(FMAP_28_36);
			MULT_37(27)<=signed(DIN_37_7)*signed(FMAP_28_37);
			MULT_38(27)<=signed(DIN_38_7)*signed(FMAP_28_38);
			MULT_39(27)<=signed(DIN_39_7)*signed(FMAP_28_39);
			MULT_40(27)<=signed(DIN_40_7)*signed(FMAP_28_40);
			MULT_41(27)<=signed(DIN_41_7)*signed(FMAP_28_41);
			MULT_42(27)<=signed(DIN_42_7)*signed(FMAP_28_42);
			MULT_43(27)<=signed(DIN_43_7)*signed(FMAP_28_43);
			MULT_44(27)<=signed(DIN_44_7)*signed(FMAP_28_44);
			MULT_45(27)<=signed(DIN_45_7)*signed(FMAP_28_45);
			MULT_46(27)<=signed(DIN_46_7)*signed(FMAP_28_46);
			MULT_47(27)<=signed(DIN_47_7)*signed(FMAP_28_47);
			MULT_48(27)<=signed(DIN_48_7)*signed(FMAP_28_48);
			MULT_49(27)<=signed(DIN_49_7)*signed(FMAP_28_49);
			MULT_50(27)<=signed(DIN_50_7)*signed(FMAP_28_50);
			MULT_51(27)<=signed(DIN_51_7)*signed(FMAP_28_51);
			MULT_52(27)<=signed(DIN_52_7)*signed(FMAP_28_52);
			MULT_53(27)<=signed(DIN_53_7)*signed(FMAP_28_53);
			MULT_54(27)<=signed(DIN_54_7)*signed(FMAP_28_54);
			MULT_55(27)<=signed(DIN_55_7)*signed(FMAP_28_55);
			MULT_56(27)<=signed(DIN_56_7)*signed(FMAP_28_56);
			MULT_57(27)<=signed(DIN_57_7)*signed(FMAP_28_57);
			MULT_58(27)<=signed(DIN_58_7)*signed(FMAP_28_58);
			MULT_59(27)<=signed(DIN_59_7)*signed(FMAP_28_59);
			MULT_60(27)<=signed(DIN_60_7)*signed(FMAP_28_60);
			MULT_61(27)<=signed(DIN_61_7)*signed(FMAP_28_61);
			MULT_62(27)<=signed(DIN_62_7)*signed(FMAP_28_62);
			MULT_63(27)<=signed(DIN_63_7)*signed(FMAP_28_63);
			MULT_64(27)<=signed(DIN_64_7)*signed(FMAP_28_64);
			MULT_65(27)<=signed(DIN_65_7)*signed(FMAP_28_65);
			MULT_66(27)<=signed(DIN_66_7)*signed(FMAP_28_66);
			MULT_67(27)<=signed(DIN_67_7)*signed(FMAP_28_67);
			MULT_68(27)<=signed(DIN_68_7)*signed(FMAP_28_68);
			MULT_69(27)<=signed(DIN_69_7)*signed(FMAP_28_69);
			MULT_70(27)<=signed(DIN_70_7)*signed(FMAP_28_70);
			MULT_71(27)<=signed(DIN_71_7)*signed(FMAP_28_71);
			MULT_72(27)<=signed(DIN_72_7)*signed(FMAP_28_72);
			MULT_73(27)<=signed(DIN_73_7)*signed(FMAP_28_73);
			MULT_74(27)<=signed(DIN_74_7)*signed(FMAP_28_74);
			MULT_75(27)<=signed(DIN_75_7)*signed(FMAP_28_75);
			MULT_76(27)<=signed(DIN_76_7)*signed(FMAP_28_76);
			MULT_77(27)<=signed(DIN_77_7)*signed(FMAP_28_77);
			MULT_78(27)<=signed(DIN_78_7)*signed(FMAP_28_78);
			MULT_79(27)<=signed(DIN_79_7)*signed(FMAP_28_79);
			MULT_80(27)<=signed(DIN_80_7)*signed(FMAP_28_80);
			MULT_81(27)<=signed(DIN_81_7)*signed(FMAP_28_81);
			MULT_82(27)<=signed(DIN_82_7)*signed(FMAP_28_82);
			MULT_83(27)<=signed(DIN_83_7)*signed(FMAP_28_83);
			MULT_84(27)<=signed(DIN_84_7)*signed(FMAP_28_84);
			MULT_85(27)<=signed(DIN_85_7)*signed(FMAP_28_85);
			MULT_86(27)<=signed(DIN_86_7)*signed(FMAP_28_86);
			MULT_87(27)<=signed(DIN_87_7)*signed(FMAP_28_87);
			MULT_88(27)<=signed(DIN_88_7)*signed(FMAP_28_88);
			MULT_89(27)<=signed(DIN_89_7)*signed(FMAP_28_89);
			MULT_90(27)<=signed(DIN_90_7)*signed(FMAP_28_90);
			MULT_91(27)<=signed(DIN_91_7)*signed(FMAP_28_91);
			MULT_92(27)<=signed(DIN_92_7)*signed(FMAP_28_92);
			MULT_93(27)<=signed(DIN_93_7)*signed(FMAP_28_93);
			MULT_94(27)<=signed(DIN_94_7)*signed(FMAP_28_94);
			MULT_95(27)<=signed(DIN_95_7)*signed(FMAP_28_95);
			MULT_96(27)<=signed(DIN_96_7)*signed(FMAP_28_96);
			MULT_97(27)<=signed(DIN_97_7)*signed(FMAP_28_97);
			MULT_98(27)<=signed(DIN_98_7)*signed(FMAP_28_98);
			MULT_99(27)<=signed(DIN_99_7)*signed(FMAP_28_99);
			MULT_100(27)<=signed(DIN_100_7)*signed(FMAP_28_100);
			MULT_101(27)<=signed(DIN_101_7)*signed(FMAP_28_101);
			MULT_102(27)<=signed(DIN_102_7)*signed(FMAP_28_102);
			MULT_103(27)<=signed(DIN_103_7)*signed(FMAP_28_103);
			MULT_104(27)<=signed(DIN_104_7)*signed(FMAP_28_104);
			MULT_105(27)<=signed(DIN_105_7)*signed(FMAP_28_105);
			MULT_106(27)<=signed(DIN_106_7)*signed(FMAP_28_106);
			MULT_107(27)<=signed(DIN_107_7)*signed(FMAP_28_107);
			MULT_108(27)<=signed(DIN_108_7)*signed(FMAP_28_108);
			MULT_109(27)<=signed(DIN_109_7)*signed(FMAP_28_109);
			MULT_110(27)<=signed(DIN_110_7)*signed(FMAP_28_110);
			MULT_111(27)<=signed(DIN_111_7)*signed(FMAP_28_111);
			MULT_112(27)<=signed(DIN_112_7)*signed(FMAP_28_112);
			MULT_113(27)<=signed(DIN_113_7)*signed(FMAP_28_113);
			MULT_114(27)<=signed(DIN_114_7)*signed(FMAP_28_114);
			MULT_115(27)<=signed(DIN_115_7)*signed(FMAP_28_115);
			MULT_116(27)<=signed(DIN_116_7)*signed(FMAP_28_116);
			MULT_117(27)<=signed(DIN_117_7)*signed(FMAP_28_117);
			MULT_118(27)<=signed(DIN_118_7)*signed(FMAP_28_118);
			MULT_119(27)<=signed(DIN_119_7)*signed(FMAP_28_119);
			MULT_120(27)<=signed(DIN_120_7)*signed(FMAP_28_120);

			MULT_1(28)<=signed(DIN_1_7)*signed(FMAP_29_1);
			MULT_2(28)<=signed(DIN_2_7)*signed(FMAP_29_2);
			MULT_3(28)<=signed(DIN_3_7)*signed(FMAP_29_3);
			MULT_4(28)<=signed(DIN_4_7)*signed(FMAP_29_4);
			MULT_5(28)<=signed(DIN_5_7)*signed(FMAP_29_5);
			MULT_6(28)<=signed(DIN_6_7)*signed(FMAP_29_6);
			MULT_7(28)<=signed(DIN_7_7)*signed(FMAP_29_7);
			MULT_8(28)<=signed(DIN_8_7)*signed(FMAP_29_8);
			MULT_9(28)<=signed(DIN_9_7)*signed(FMAP_29_9);
			MULT_10(28)<=signed(DIN_10_7)*signed(FMAP_29_10);
			MULT_11(28)<=signed(DIN_11_7)*signed(FMAP_29_11);
			MULT_12(28)<=signed(DIN_12_7)*signed(FMAP_29_12);
			MULT_13(28)<=signed(DIN_13_7)*signed(FMAP_29_13);
			MULT_14(28)<=signed(DIN_14_7)*signed(FMAP_29_14);
			MULT_15(28)<=signed(DIN_15_7)*signed(FMAP_29_15);
			MULT_16(28)<=signed(DIN_16_7)*signed(FMAP_29_16);
			MULT_17(28)<=signed(DIN_17_7)*signed(FMAP_29_17);
			MULT_18(28)<=signed(DIN_18_7)*signed(FMAP_29_18);
			MULT_19(28)<=signed(DIN_19_7)*signed(FMAP_29_19);
			MULT_20(28)<=signed(DIN_20_7)*signed(FMAP_29_20);
			MULT_21(28)<=signed(DIN_21_7)*signed(FMAP_29_21);
			MULT_22(28)<=signed(DIN_22_7)*signed(FMAP_29_22);
			MULT_23(28)<=signed(DIN_23_7)*signed(FMAP_29_23);
			MULT_24(28)<=signed(DIN_24_7)*signed(FMAP_29_24);
			MULT_25(28)<=signed(DIN_25_7)*signed(FMAP_29_25);
			MULT_26(28)<=signed(DIN_26_7)*signed(FMAP_29_26);
			MULT_27(28)<=signed(DIN_27_7)*signed(FMAP_29_27);
			MULT_28(28)<=signed(DIN_28_7)*signed(FMAP_29_28);
			MULT_29(28)<=signed(DIN_29_7)*signed(FMAP_29_29);
			MULT_30(28)<=signed(DIN_30_7)*signed(FMAP_29_30);
			MULT_31(28)<=signed(DIN_31_7)*signed(FMAP_29_31);
			MULT_32(28)<=signed(DIN_32_7)*signed(FMAP_29_32);
			MULT_33(28)<=signed(DIN_33_7)*signed(FMAP_29_33);
			MULT_34(28)<=signed(DIN_34_7)*signed(FMAP_29_34);
			MULT_35(28)<=signed(DIN_35_7)*signed(FMAP_29_35);
			MULT_36(28)<=signed(DIN_36_7)*signed(FMAP_29_36);
			MULT_37(28)<=signed(DIN_37_7)*signed(FMAP_29_37);
			MULT_38(28)<=signed(DIN_38_7)*signed(FMAP_29_38);
			MULT_39(28)<=signed(DIN_39_7)*signed(FMAP_29_39);
			MULT_40(28)<=signed(DIN_40_7)*signed(FMAP_29_40);
			MULT_41(28)<=signed(DIN_41_7)*signed(FMAP_29_41);
			MULT_42(28)<=signed(DIN_42_7)*signed(FMAP_29_42);
			MULT_43(28)<=signed(DIN_43_7)*signed(FMAP_29_43);
			MULT_44(28)<=signed(DIN_44_7)*signed(FMAP_29_44);
			MULT_45(28)<=signed(DIN_45_7)*signed(FMAP_29_45);
			MULT_46(28)<=signed(DIN_46_7)*signed(FMAP_29_46);
			MULT_47(28)<=signed(DIN_47_7)*signed(FMAP_29_47);
			MULT_48(28)<=signed(DIN_48_7)*signed(FMAP_29_48);
			MULT_49(28)<=signed(DIN_49_7)*signed(FMAP_29_49);
			MULT_50(28)<=signed(DIN_50_7)*signed(FMAP_29_50);
			MULT_51(28)<=signed(DIN_51_7)*signed(FMAP_29_51);
			MULT_52(28)<=signed(DIN_52_7)*signed(FMAP_29_52);
			MULT_53(28)<=signed(DIN_53_7)*signed(FMAP_29_53);
			MULT_54(28)<=signed(DIN_54_7)*signed(FMAP_29_54);
			MULT_55(28)<=signed(DIN_55_7)*signed(FMAP_29_55);
			MULT_56(28)<=signed(DIN_56_7)*signed(FMAP_29_56);
			MULT_57(28)<=signed(DIN_57_7)*signed(FMAP_29_57);
			MULT_58(28)<=signed(DIN_58_7)*signed(FMAP_29_58);
			MULT_59(28)<=signed(DIN_59_7)*signed(FMAP_29_59);
			MULT_60(28)<=signed(DIN_60_7)*signed(FMAP_29_60);
			MULT_61(28)<=signed(DIN_61_7)*signed(FMAP_29_61);
			MULT_62(28)<=signed(DIN_62_7)*signed(FMAP_29_62);
			MULT_63(28)<=signed(DIN_63_7)*signed(FMAP_29_63);
			MULT_64(28)<=signed(DIN_64_7)*signed(FMAP_29_64);
			MULT_65(28)<=signed(DIN_65_7)*signed(FMAP_29_65);
			MULT_66(28)<=signed(DIN_66_7)*signed(FMAP_29_66);
			MULT_67(28)<=signed(DIN_67_7)*signed(FMAP_29_67);
			MULT_68(28)<=signed(DIN_68_7)*signed(FMAP_29_68);
			MULT_69(28)<=signed(DIN_69_7)*signed(FMAP_29_69);
			MULT_70(28)<=signed(DIN_70_7)*signed(FMAP_29_70);
			MULT_71(28)<=signed(DIN_71_7)*signed(FMAP_29_71);
			MULT_72(28)<=signed(DIN_72_7)*signed(FMAP_29_72);
			MULT_73(28)<=signed(DIN_73_7)*signed(FMAP_29_73);
			MULT_74(28)<=signed(DIN_74_7)*signed(FMAP_29_74);
			MULT_75(28)<=signed(DIN_75_7)*signed(FMAP_29_75);
			MULT_76(28)<=signed(DIN_76_7)*signed(FMAP_29_76);
			MULT_77(28)<=signed(DIN_77_7)*signed(FMAP_29_77);
			MULT_78(28)<=signed(DIN_78_7)*signed(FMAP_29_78);
			MULT_79(28)<=signed(DIN_79_7)*signed(FMAP_29_79);
			MULT_80(28)<=signed(DIN_80_7)*signed(FMAP_29_80);
			MULT_81(28)<=signed(DIN_81_7)*signed(FMAP_29_81);
			MULT_82(28)<=signed(DIN_82_7)*signed(FMAP_29_82);
			MULT_83(28)<=signed(DIN_83_7)*signed(FMAP_29_83);
			MULT_84(28)<=signed(DIN_84_7)*signed(FMAP_29_84);
			MULT_85(28)<=signed(DIN_85_7)*signed(FMAP_29_85);
			MULT_86(28)<=signed(DIN_86_7)*signed(FMAP_29_86);
			MULT_87(28)<=signed(DIN_87_7)*signed(FMAP_29_87);
			MULT_88(28)<=signed(DIN_88_7)*signed(FMAP_29_88);
			MULT_89(28)<=signed(DIN_89_7)*signed(FMAP_29_89);
			MULT_90(28)<=signed(DIN_90_7)*signed(FMAP_29_90);
			MULT_91(28)<=signed(DIN_91_7)*signed(FMAP_29_91);
			MULT_92(28)<=signed(DIN_92_7)*signed(FMAP_29_92);
			MULT_93(28)<=signed(DIN_93_7)*signed(FMAP_29_93);
			MULT_94(28)<=signed(DIN_94_7)*signed(FMAP_29_94);
			MULT_95(28)<=signed(DIN_95_7)*signed(FMAP_29_95);
			MULT_96(28)<=signed(DIN_96_7)*signed(FMAP_29_96);
			MULT_97(28)<=signed(DIN_97_7)*signed(FMAP_29_97);
			MULT_98(28)<=signed(DIN_98_7)*signed(FMAP_29_98);
			MULT_99(28)<=signed(DIN_99_7)*signed(FMAP_29_99);
			MULT_100(28)<=signed(DIN_100_7)*signed(FMAP_29_100);
			MULT_101(28)<=signed(DIN_101_7)*signed(FMAP_29_101);
			MULT_102(28)<=signed(DIN_102_7)*signed(FMAP_29_102);
			MULT_103(28)<=signed(DIN_103_7)*signed(FMAP_29_103);
			MULT_104(28)<=signed(DIN_104_7)*signed(FMAP_29_104);
			MULT_105(28)<=signed(DIN_105_7)*signed(FMAP_29_105);
			MULT_106(28)<=signed(DIN_106_7)*signed(FMAP_29_106);
			MULT_107(28)<=signed(DIN_107_7)*signed(FMAP_29_107);
			MULT_108(28)<=signed(DIN_108_7)*signed(FMAP_29_108);
			MULT_109(28)<=signed(DIN_109_7)*signed(FMAP_29_109);
			MULT_110(28)<=signed(DIN_110_7)*signed(FMAP_29_110);
			MULT_111(28)<=signed(DIN_111_7)*signed(FMAP_29_111);
			MULT_112(28)<=signed(DIN_112_7)*signed(FMAP_29_112);
			MULT_113(28)<=signed(DIN_113_7)*signed(FMAP_29_113);
			MULT_114(28)<=signed(DIN_114_7)*signed(FMAP_29_114);
			MULT_115(28)<=signed(DIN_115_7)*signed(FMAP_29_115);
			MULT_116(28)<=signed(DIN_116_7)*signed(FMAP_29_116);
			MULT_117(28)<=signed(DIN_117_7)*signed(FMAP_29_117);
			MULT_118(28)<=signed(DIN_118_7)*signed(FMAP_29_118);
			MULT_119(28)<=signed(DIN_119_7)*signed(FMAP_29_119);
			MULT_120(28)<=signed(DIN_120_7)*signed(FMAP_29_120);

			MULT_1(29)<=signed(DIN_1_7)*signed(FMAP_30_1);
			MULT_2(29)<=signed(DIN_2_7)*signed(FMAP_30_2);
			MULT_3(29)<=signed(DIN_3_7)*signed(FMAP_30_3);
			MULT_4(29)<=signed(DIN_4_7)*signed(FMAP_30_4);
			MULT_5(29)<=signed(DIN_5_7)*signed(FMAP_30_5);
			MULT_6(29)<=signed(DIN_6_7)*signed(FMAP_30_6);
			MULT_7(29)<=signed(DIN_7_7)*signed(FMAP_30_7);
			MULT_8(29)<=signed(DIN_8_7)*signed(FMAP_30_8);
			MULT_9(29)<=signed(DIN_9_7)*signed(FMAP_30_9);
			MULT_10(29)<=signed(DIN_10_7)*signed(FMAP_30_10);
			MULT_11(29)<=signed(DIN_11_7)*signed(FMAP_30_11);
			MULT_12(29)<=signed(DIN_12_7)*signed(FMAP_30_12);
			MULT_13(29)<=signed(DIN_13_7)*signed(FMAP_30_13);
			MULT_14(29)<=signed(DIN_14_7)*signed(FMAP_30_14);
			MULT_15(29)<=signed(DIN_15_7)*signed(FMAP_30_15);
			MULT_16(29)<=signed(DIN_16_7)*signed(FMAP_30_16);
			MULT_17(29)<=signed(DIN_17_7)*signed(FMAP_30_17);
			MULT_18(29)<=signed(DIN_18_7)*signed(FMAP_30_18);
			MULT_19(29)<=signed(DIN_19_7)*signed(FMAP_30_19);
			MULT_20(29)<=signed(DIN_20_7)*signed(FMAP_30_20);
			MULT_21(29)<=signed(DIN_21_7)*signed(FMAP_30_21);
			MULT_22(29)<=signed(DIN_22_7)*signed(FMAP_30_22);
			MULT_23(29)<=signed(DIN_23_7)*signed(FMAP_30_23);
			MULT_24(29)<=signed(DIN_24_7)*signed(FMAP_30_24);
			MULT_25(29)<=signed(DIN_25_7)*signed(FMAP_30_25);
			MULT_26(29)<=signed(DIN_26_7)*signed(FMAP_30_26);
			MULT_27(29)<=signed(DIN_27_7)*signed(FMAP_30_27);
			MULT_28(29)<=signed(DIN_28_7)*signed(FMAP_30_28);
			MULT_29(29)<=signed(DIN_29_7)*signed(FMAP_30_29);
			MULT_30(29)<=signed(DIN_30_7)*signed(FMAP_30_30);
			MULT_31(29)<=signed(DIN_31_7)*signed(FMAP_30_31);
			MULT_32(29)<=signed(DIN_32_7)*signed(FMAP_30_32);
			MULT_33(29)<=signed(DIN_33_7)*signed(FMAP_30_33);
			MULT_34(29)<=signed(DIN_34_7)*signed(FMAP_30_34);
			MULT_35(29)<=signed(DIN_35_7)*signed(FMAP_30_35);
			MULT_36(29)<=signed(DIN_36_7)*signed(FMAP_30_36);
			MULT_37(29)<=signed(DIN_37_7)*signed(FMAP_30_37);
			MULT_38(29)<=signed(DIN_38_7)*signed(FMAP_30_38);
			MULT_39(29)<=signed(DIN_39_7)*signed(FMAP_30_39);
			MULT_40(29)<=signed(DIN_40_7)*signed(FMAP_30_40);
			MULT_41(29)<=signed(DIN_41_7)*signed(FMAP_30_41);
			MULT_42(29)<=signed(DIN_42_7)*signed(FMAP_30_42);
			MULT_43(29)<=signed(DIN_43_7)*signed(FMAP_30_43);
			MULT_44(29)<=signed(DIN_44_7)*signed(FMAP_30_44);
			MULT_45(29)<=signed(DIN_45_7)*signed(FMAP_30_45);
			MULT_46(29)<=signed(DIN_46_7)*signed(FMAP_30_46);
			MULT_47(29)<=signed(DIN_47_7)*signed(FMAP_30_47);
			MULT_48(29)<=signed(DIN_48_7)*signed(FMAP_30_48);
			MULT_49(29)<=signed(DIN_49_7)*signed(FMAP_30_49);
			MULT_50(29)<=signed(DIN_50_7)*signed(FMAP_30_50);
			MULT_51(29)<=signed(DIN_51_7)*signed(FMAP_30_51);
			MULT_52(29)<=signed(DIN_52_7)*signed(FMAP_30_52);
			MULT_53(29)<=signed(DIN_53_7)*signed(FMAP_30_53);
			MULT_54(29)<=signed(DIN_54_7)*signed(FMAP_30_54);
			MULT_55(29)<=signed(DIN_55_7)*signed(FMAP_30_55);
			MULT_56(29)<=signed(DIN_56_7)*signed(FMAP_30_56);
			MULT_57(29)<=signed(DIN_57_7)*signed(FMAP_30_57);
			MULT_58(29)<=signed(DIN_58_7)*signed(FMAP_30_58);
			MULT_59(29)<=signed(DIN_59_7)*signed(FMAP_30_59);
			MULT_60(29)<=signed(DIN_60_7)*signed(FMAP_30_60);
			MULT_61(29)<=signed(DIN_61_7)*signed(FMAP_30_61);
			MULT_62(29)<=signed(DIN_62_7)*signed(FMAP_30_62);
			MULT_63(29)<=signed(DIN_63_7)*signed(FMAP_30_63);
			MULT_64(29)<=signed(DIN_64_7)*signed(FMAP_30_64);
			MULT_65(29)<=signed(DIN_65_7)*signed(FMAP_30_65);
			MULT_66(29)<=signed(DIN_66_7)*signed(FMAP_30_66);
			MULT_67(29)<=signed(DIN_67_7)*signed(FMAP_30_67);
			MULT_68(29)<=signed(DIN_68_7)*signed(FMAP_30_68);
			MULT_69(29)<=signed(DIN_69_7)*signed(FMAP_30_69);
			MULT_70(29)<=signed(DIN_70_7)*signed(FMAP_30_70);
			MULT_71(29)<=signed(DIN_71_7)*signed(FMAP_30_71);
			MULT_72(29)<=signed(DIN_72_7)*signed(FMAP_30_72);
			MULT_73(29)<=signed(DIN_73_7)*signed(FMAP_30_73);
			MULT_74(29)<=signed(DIN_74_7)*signed(FMAP_30_74);
			MULT_75(29)<=signed(DIN_75_7)*signed(FMAP_30_75);
			MULT_76(29)<=signed(DIN_76_7)*signed(FMAP_30_76);
			MULT_77(29)<=signed(DIN_77_7)*signed(FMAP_30_77);
			MULT_78(29)<=signed(DIN_78_7)*signed(FMAP_30_78);
			MULT_79(29)<=signed(DIN_79_7)*signed(FMAP_30_79);
			MULT_80(29)<=signed(DIN_80_7)*signed(FMAP_30_80);
			MULT_81(29)<=signed(DIN_81_7)*signed(FMAP_30_81);
			MULT_82(29)<=signed(DIN_82_7)*signed(FMAP_30_82);
			MULT_83(29)<=signed(DIN_83_7)*signed(FMAP_30_83);
			MULT_84(29)<=signed(DIN_84_7)*signed(FMAP_30_84);
			MULT_85(29)<=signed(DIN_85_7)*signed(FMAP_30_85);
			MULT_86(29)<=signed(DIN_86_7)*signed(FMAP_30_86);
			MULT_87(29)<=signed(DIN_87_7)*signed(FMAP_30_87);
			MULT_88(29)<=signed(DIN_88_7)*signed(FMAP_30_88);
			MULT_89(29)<=signed(DIN_89_7)*signed(FMAP_30_89);
			MULT_90(29)<=signed(DIN_90_7)*signed(FMAP_30_90);
			MULT_91(29)<=signed(DIN_91_7)*signed(FMAP_30_91);
			MULT_92(29)<=signed(DIN_92_7)*signed(FMAP_30_92);
			MULT_93(29)<=signed(DIN_93_7)*signed(FMAP_30_93);
			MULT_94(29)<=signed(DIN_94_7)*signed(FMAP_30_94);
			MULT_95(29)<=signed(DIN_95_7)*signed(FMAP_30_95);
			MULT_96(29)<=signed(DIN_96_7)*signed(FMAP_30_96);
			MULT_97(29)<=signed(DIN_97_7)*signed(FMAP_30_97);
			MULT_98(29)<=signed(DIN_98_7)*signed(FMAP_30_98);
			MULT_99(29)<=signed(DIN_99_7)*signed(FMAP_30_99);
			MULT_100(29)<=signed(DIN_100_7)*signed(FMAP_30_100);
			MULT_101(29)<=signed(DIN_101_7)*signed(FMAP_30_101);
			MULT_102(29)<=signed(DIN_102_7)*signed(FMAP_30_102);
			MULT_103(29)<=signed(DIN_103_7)*signed(FMAP_30_103);
			MULT_104(29)<=signed(DIN_104_7)*signed(FMAP_30_104);
			MULT_105(29)<=signed(DIN_105_7)*signed(FMAP_30_105);
			MULT_106(29)<=signed(DIN_106_7)*signed(FMAP_30_106);
			MULT_107(29)<=signed(DIN_107_7)*signed(FMAP_30_107);
			MULT_108(29)<=signed(DIN_108_7)*signed(FMAP_30_108);
			MULT_109(29)<=signed(DIN_109_7)*signed(FMAP_30_109);
			MULT_110(29)<=signed(DIN_110_7)*signed(FMAP_30_110);
			MULT_111(29)<=signed(DIN_111_7)*signed(FMAP_30_111);
			MULT_112(29)<=signed(DIN_112_7)*signed(FMAP_30_112);
			MULT_113(29)<=signed(DIN_113_7)*signed(FMAP_30_113);
			MULT_114(29)<=signed(DIN_114_7)*signed(FMAP_30_114);
			MULT_115(29)<=signed(DIN_115_7)*signed(FMAP_30_115);
			MULT_116(29)<=signed(DIN_116_7)*signed(FMAP_30_116);
			MULT_117(29)<=signed(DIN_117_7)*signed(FMAP_30_117);
			MULT_118(29)<=signed(DIN_118_7)*signed(FMAP_30_118);
			MULT_119(29)<=signed(DIN_119_7)*signed(FMAP_30_119);
			MULT_120(29)<=signed(DIN_120_7)*signed(FMAP_30_120);

			MULT_1(30)<=signed(DIN_1_7)*signed(FMAP_31_1);
			MULT_2(30)<=signed(DIN_2_7)*signed(FMAP_31_2);
			MULT_3(30)<=signed(DIN_3_7)*signed(FMAP_31_3);
			MULT_4(30)<=signed(DIN_4_7)*signed(FMAP_31_4);
			MULT_5(30)<=signed(DIN_5_7)*signed(FMAP_31_5);
			MULT_6(30)<=signed(DIN_6_7)*signed(FMAP_31_6);
			MULT_7(30)<=signed(DIN_7_7)*signed(FMAP_31_7);
			MULT_8(30)<=signed(DIN_8_7)*signed(FMAP_31_8);
			MULT_9(30)<=signed(DIN_9_7)*signed(FMAP_31_9);
			MULT_10(30)<=signed(DIN_10_7)*signed(FMAP_31_10);
			MULT_11(30)<=signed(DIN_11_7)*signed(FMAP_31_11);
			MULT_12(30)<=signed(DIN_12_7)*signed(FMAP_31_12);
			MULT_13(30)<=signed(DIN_13_7)*signed(FMAP_31_13);
			MULT_14(30)<=signed(DIN_14_7)*signed(FMAP_31_14);
			MULT_15(30)<=signed(DIN_15_7)*signed(FMAP_31_15);
			MULT_16(30)<=signed(DIN_16_7)*signed(FMAP_31_16);
			MULT_17(30)<=signed(DIN_17_7)*signed(FMAP_31_17);
			MULT_18(30)<=signed(DIN_18_7)*signed(FMAP_31_18);
			MULT_19(30)<=signed(DIN_19_7)*signed(FMAP_31_19);
			MULT_20(30)<=signed(DIN_20_7)*signed(FMAP_31_20);
			MULT_21(30)<=signed(DIN_21_7)*signed(FMAP_31_21);
			MULT_22(30)<=signed(DIN_22_7)*signed(FMAP_31_22);
			MULT_23(30)<=signed(DIN_23_7)*signed(FMAP_31_23);
			MULT_24(30)<=signed(DIN_24_7)*signed(FMAP_31_24);
			MULT_25(30)<=signed(DIN_25_7)*signed(FMAP_31_25);
			MULT_26(30)<=signed(DIN_26_7)*signed(FMAP_31_26);
			MULT_27(30)<=signed(DIN_27_7)*signed(FMAP_31_27);
			MULT_28(30)<=signed(DIN_28_7)*signed(FMAP_31_28);
			MULT_29(30)<=signed(DIN_29_7)*signed(FMAP_31_29);
			MULT_30(30)<=signed(DIN_30_7)*signed(FMAP_31_30);
			MULT_31(30)<=signed(DIN_31_7)*signed(FMAP_31_31);
			MULT_32(30)<=signed(DIN_32_7)*signed(FMAP_31_32);
			MULT_33(30)<=signed(DIN_33_7)*signed(FMAP_31_33);
			MULT_34(30)<=signed(DIN_34_7)*signed(FMAP_31_34);
			MULT_35(30)<=signed(DIN_35_7)*signed(FMAP_31_35);
			MULT_36(30)<=signed(DIN_36_7)*signed(FMAP_31_36);
			MULT_37(30)<=signed(DIN_37_7)*signed(FMAP_31_37);
			MULT_38(30)<=signed(DIN_38_7)*signed(FMAP_31_38);
			MULT_39(30)<=signed(DIN_39_7)*signed(FMAP_31_39);
			MULT_40(30)<=signed(DIN_40_7)*signed(FMAP_31_40);
			MULT_41(30)<=signed(DIN_41_7)*signed(FMAP_31_41);
			MULT_42(30)<=signed(DIN_42_7)*signed(FMAP_31_42);
			MULT_43(30)<=signed(DIN_43_7)*signed(FMAP_31_43);
			MULT_44(30)<=signed(DIN_44_7)*signed(FMAP_31_44);
			MULT_45(30)<=signed(DIN_45_7)*signed(FMAP_31_45);
			MULT_46(30)<=signed(DIN_46_7)*signed(FMAP_31_46);
			MULT_47(30)<=signed(DIN_47_7)*signed(FMAP_31_47);
			MULT_48(30)<=signed(DIN_48_7)*signed(FMAP_31_48);
			MULT_49(30)<=signed(DIN_49_7)*signed(FMAP_31_49);
			MULT_50(30)<=signed(DIN_50_7)*signed(FMAP_31_50);
			MULT_51(30)<=signed(DIN_51_7)*signed(FMAP_31_51);
			MULT_52(30)<=signed(DIN_52_7)*signed(FMAP_31_52);
			MULT_53(30)<=signed(DIN_53_7)*signed(FMAP_31_53);
			MULT_54(30)<=signed(DIN_54_7)*signed(FMAP_31_54);
			MULT_55(30)<=signed(DIN_55_7)*signed(FMAP_31_55);
			MULT_56(30)<=signed(DIN_56_7)*signed(FMAP_31_56);
			MULT_57(30)<=signed(DIN_57_7)*signed(FMAP_31_57);
			MULT_58(30)<=signed(DIN_58_7)*signed(FMAP_31_58);
			MULT_59(30)<=signed(DIN_59_7)*signed(FMAP_31_59);
			MULT_60(30)<=signed(DIN_60_7)*signed(FMAP_31_60);
			MULT_61(30)<=signed(DIN_61_7)*signed(FMAP_31_61);
			MULT_62(30)<=signed(DIN_62_7)*signed(FMAP_31_62);
			MULT_63(30)<=signed(DIN_63_7)*signed(FMAP_31_63);
			MULT_64(30)<=signed(DIN_64_7)*signed(FMAP_31_64);
			MULT_65(30)<=signed(DIN_65_7)*signed(FMAP_31_65);
			MULT_66(30)<=signed(DIN_66_7)*signed(FMAP_31_66);
			MULT_67(30)<=signed(DIN_67_7)*signed(FMAP_31_67);
			MULT_68(30)<=signed(DIN_68_7)*signed(FMAP_31_68);
			MULT_69(30)<=signed(DIN_69_7)*signed(FMAP_31_69);
			MULT_70(30)<=signed(DIN_70_7)*signed(FMAP_31_70);
			MULT_71(30)<=signed(DIN_71_7)*signed(FMAP_31_71);
			MULT_72(30)<=signed(DIN_72_7)*signed(FMAP_31_72);
			MULT_73(30)<=signed(DIN_73_7)*signed(FMAP_31_73);
			MULT_74(30)<=signed(DIN_74_7)*signed(FMAP_31_74);
			MULT_75(30)<=signed(DIN_75_7)*signed(FMAP_31_75);
			MULT_76(30)<=signed(DIN_76_7)*signed(FMAP_31_76);
			MULT_77(30)<=signed(DIN_77_7)*signed(FMAP_31_77);
			MULT_78(30)<=signed(DIN_78_7)*signed(FMAP_31_78);
			MULT_79(30)<=signed(DIN_79_7)*signed(FMAP_31_79);
			MULT_80(30)<=signed(DIN_80_7)*signed(FMAP_31_80);
			MULT_81(30)<=signed(DIN_81_7)*signed(FMAP_31_81);
			MULT_82(30)<=signed(DIN_82_7)*signed(FMAP_31_82);
			MULT_83(30)<=signed(DIN_83_7)*signed(FMAP_31_83);
			MULT_84(30)<=signed(DIN_84_7)*signed(FMAP_31_84);
			MULT_85(30)<=signed(DIN_85_7)*signed(FMAP_31_85);
			MULT_86(30)<=signed(DIN_86_7)*signed(FMAP_31_86);
			MULT_87(30)<=signed(DIN_87_7)*signed(FMAP_31_87);
			MULT_88(30)<=signed(DIN_88_7)*signed(FMAP_31_88);
			MULT_89(30)<=signed(DIN_89_7)*signed(FMAP_31_89);
			MULT_90(30)<=signed(DIN_90_7)*signed(FMAP_31_90);
			MULT_91(30)<=signed(DIN_91_7)*signed(FMAP_31_91);
			MULT_92(30)<=signed(DIN_92_7)*signed(FMAP_31_92);
			MULT_93(30)<=signed(DIN_93_7)*signed(FMAP_31_93);
			MULT_94(30)<=signed(DIN_94_7)*signed(FMAP_31_94);
			MULT_95(30)<=signed(DIN_95_7)*signed(FMAP_31_95);
			MULT_96(30)<=signed(DIN_96_7)*signed(FMAP_31_96);
			MULT_97(30)<=signed(DIN_97_7)*signed(FMAP_31_97);
			MULT_98(30)<=signed(DIN_98_7)*signed(FMAP_31_98);
			MULT_99(30)<=signed(DIN_99_7)*signed(FMAP_31_99);
			MULT_100(30)<=signed(DIN_100_7)*signed(FMAP_31_100);
			MULT_101(30)<=signed(DIN_101_7)*signed(FMAP_31_101);
			MULT_102(30)<=signed(DIN_102_7)*signed(FMAP_31_102);
			MULT_103(30)<=signed(DIN_103_7)*signed(FMAP_31_103);
			MULT_104(30)<=signed(DIN_104_7)*signed(FMAP_31_104);
			MULT_105(30)<=signed(DIN_105_7)*signed(FMAP_31_105);
			MULT_106(30)<=signed(DIN_106_7)*signed(FMAP_31_106);
			MULT_107(30)<=signed(DIN_107_7)*signed(FMAP_31_107);
			MULT_108(30)<=signed(DIN_108_7)*signed(FMAP_31_108);
			MULT_109(30)<=signed(DIN_109_7)*signed(FMAP_31_109);
			MULT_110(30)<=signed(DIN_110_7)*signed(FMAP_31_110);
			MULT_111(30)<=signed(DIN_111_7)*signed(FMAP_31_111);
			MULT_112(30)<=signed(DIN_112_7)*signed(FMAP_31_112);
			MULT_113(30)<=signed(DIN_113_7)*signed(FMAP_31_113);
			MULT_114(30)<=signed(DIN_114_7)*signed(FMAP_31_114);
			MULT_115(30)<=signed(DIN_115_7)*signed(FMAP_31_115);
			MULT_116(30)<=signed(DIN_116_7)*signed(FMAP_31_116);
			MULT_117(30)<=signed(DIN_117_7)*signed(FMAP_31_117);
			MULT_118(30)<=signed(DIN_118_7)*signed(FMAP_31_118);
			MULT_119(30)<=signed(DIN_119_7)*signed(FMAP_31_119);
			MULT_120(30)<=signed(DIN_120_7)*signed(FMAP_31_120);

			MULT_1(31)<=signed(DIN_1_7)*signed(FMAP_32_1);
			MULT_2(31)<=signed(DIN_2_7)*signed(FMAP_32_2);
			MULT_3(31)<=signed(DIN_3_7)*signed(FMAP_32_3);
			MULT_4(31)<=signed(DIN_4_7)*signed(FMAP_32_4);
			MULT_5(31)<=signed(DIN_5_7)*signed(FMAP_32_5);
			MULT_6(31)<=signed(DIN_6_7)*signed(FMAP_32_6);
			MULT_7(31)<=signed(DIN_7_7)*signed(FMAP_32_7);
			MULT_8(31)<=signed(DIN_8_7)*signed(FMAP_32_8);
			MULT_9(31)<=signed(DIN_9_7)*signed(FMAP_32_9);
			MULT_10(31)<=signed(DIN_10_7)*signed(FMAP_32_10);
			MULT_11(31)<=signed(DIN_11_7)*signed(FMAP_32_11);
			MULT_12(31)<=signed(DIN_12_7)*signed(FMAP_32_12);
			MULT_13(31)<=signed(DIN_13_7)*signed(FMAP_32_13);
			MULT_14(31)<=signed(DIN_14_7)*signed(FMAP_32_14);
			MULT_15(31)<=signed(DIN_15_7)*signed(FMAP_32_15);
			MULT_16(31)<=signed(DIN_16_7)*signed(FMAP_32_16);
			MULT_17(31)<=signed(DIN_17_7)*signed(FMAP_32_17);
			MULT_18(31)<=signed(DIN_18_7)*signed(FMAP_32_18);
			MULT_19(31)<=signed(DIN_19_7)*signed(FMAP_32_19);
			MULT_20(31)<=signed(DIN_20_7)*signed(FMAP_32_20);
			MULT_21(31)<=signed(DIN_21_7)*signed(FMAP_32_21);
			MULT_22(31)<=signed(DIN_22_7)*signed(FMAP_32_22);
			MULT_23(31)<=signed(DIN_23_7)*signed(FMAP_32_23);
			MULT_24(31)<=signed(DIN_24_7)*signed(FMAP_32_24);
			MULT_25(31)<=signed(DIN_25_7)*signed(FMAP_32_25);
			MULT_26(31)<=signed(DIN_26_7)*signed(FMAP_32_26);
			MULT_27(31)<=signed(DIN_27_7)*signed(FMAP_32_27);
			MULT_28(31)<=signed(DIN_28_7)*signed(FMAP_32_28);
			MULT_29(31)<=signed(DIN_29_7)*signed(FMAP_32_29);
			MULT_30(31)<=signed(DIN_30_7)*signed(FMAP_32_30);
			MULT_31(31)<=signed(DIN_31_7)*signed(FMAP_32_31);
			MULT_32(31)<=signed(DIN_32_7)*signed(FMAP_32_32);
			MULT_33(31)<=signed(DIN_33_7)*signed(FMAP_32_33);
			MULT_34(31)<=signed(DIN_34_7)*signed(FMAP_32_34);
			MULT_35(31)<=signed(DIN_35_7)*signed(FMAP_32_35);
			MULT_36(31)<=signed(DIN_36_7)*signed(FMAP_32_36);
			MULT_37(31)<=signed(DIN_37_7)*signed(FMAP_32_37);
			MULT_38(31)<=signed(DIN_38_7)*signed(FMAP_32_38);
			MULT_39(31)<=signed(DIN_39_7)*signed(FMAP_32_39);
			MULT_40(31)<=signed(DIN_40_7)*signed(FMAP_32_40);
			MULT_41(31)<=signed(DIN_41_7)*signed(FMAP_32_41);
			MULT_42(31)<=signed(DIN_42_7)*signed(FMAP_32_42);
			MULT_43(31)<=signed(DIN_43_7)*signed(FMAP_32_43);
			MULT_44(31)<=signed(DIN_44_7)*signed(FMAP_32_44);
			MULT_45(31)<=signed(DIN_45_7)*signed(FMAP_32_45);
			MULT_46(31)<=signed(DIN_46_7)*signed(FMAP_32_46);
			MULT_47(31)<=signed(DIN_47_7)*signed(FMAP_32_47);
			MULT_48(31)<=signed(DIN_48_7)*signed(FMAP_32_48);
			MULT_49(31)<=signed(DIN_49_7)*signed(FMAP_32_49);
			MULT_50(31)<=signed(DIN_50_7)*signed(FMAP_32_50);
			MULT_51(31)<=signed(DIN_51_7)*signed(FMAP_32_51);
			MULT_52(31)<=signed(DIN_52_7)*signed(FMAP_32_52);
			MULT_53(31)<=signed(DIN_53_7)*signed(FMAP_32_53);
			MULT_54(31)<=signed(DIN_54_7)*signed(FMAP_32_54);
			MULT_55(31)<=signed(DIN_55_7)*signed(FMAP_32_55);
			MULT_56(31)<=signed(DIN_56_7)*signed(FMAP_32_56);
			MULT_57(31)<=signed(DIN_57_7)*signed(FMAP_32_57);
			MULT_58(31)<=signed(DIN_58_7)*signed(FMAP_32_58);
			MULT_59(31)<=signed(DIN_59_7)*signed(FMAP_32_59);
			MULT_60(31)<=signed(DIN_60_7)*signed(FMAP_32_60);
			MULT_61(31)<=signed(DIN_61_7)*signed(FMAP_32_61);
			MULT_62(31)<=signed(DIN_62_7)*signed(FMAP_32_62);
			MULT_63(31)<=signed(DIN_63_7)*signed(FMAP_32_63);
			MULT_64(31)<=signed(DIN_64_7)*signed(FMAP_32_64);
			MULT_65(31)<=signed(DIN_65_7)*signed(FMAP_32_65);
			MULT_66(31)<=signed(DIN_66_7)*signed(FMAP_32_66);
			MULT_67(31)<=signed(DIN_67_7)*signed(FMAP_32_67);
			MULT_68(31)<=signed(DIN_68_7)*signed(FMAP_32_68);
			MULT_69(31)<=signed(DIN_69_7)*signed(FMAP_32_69);
			MULT_70(31)<=signed(DIN_70_7)*signed(FMAP_32_70);
			MULT_71(31)<=signed(DIN_71_7)*signed(FMAP_32_71);
			MULT_72(31)<=signed(DIN_72_7)*signed(FMAP_32_72);
			MULT_73(31)<=signed(DIN_73_7)*signed(FMAP_32_73);
			MULT_74(31)<=signed(DIN_74_7)*signed(FMAP_32_74);
			MULT_75(31)<=signed(DIN_75_7)*signed(FMAP_32_75);
			MULT_76(31)<=signed(DIN_76_7)*signed(FMAP_32_76);
			MULT_77(31)<=signed(DIN_77_7)*signed(FMAP_32_77);
			MULT_78(31)<=signed(DIN_78_7)*signed(FMAP_32_78);
			MULT_79(31)<=signed(DIN_79_7)*signed(FMAP_32_79);
			MULT_80(31)<=signed(DIN_80_7)*signed(FMAP_32_80);
			MULT_81(31)<=signed(DIN_81_7)*signed(FMAP_32_81);
			MULT_82(31)<=signed(DIN_82_7)*signed(FMAP_32_82);
			MULT_83(31)<=signed(DIN_83_7)*signed(FMAP_32_83);
			MULT_84(31)<=signed(DIN_84_7)*signed(FMAP_32_84);
			MULT_85(31)<=signed(DIN_85_7)*signed(FMAP_32_85);
			MULT_86(31)<=signed(DIN_86_7)*signed(FMAP_32_86);
			MULT_87(31)<=signed(DIN_87_7)*signed(FMAP_32_87);
			MULT_88(31)<=signed(DIN_88_7)*signed(FMAP_32_88);
			MULT_89(31)<=signed(DIN_89_7)*signed(FMAP_32_89);
			MULT_90(31)<=signed(DIN_90_7)*signed(FMAP_32_90);
			MULT_91(31)<=signed(DIN_91_7)*signed(FMAP_32_91);
			MULT_92(31)<=signed(DIN_92_7)*signed(FMAP_32_92);
			MULT_93(31)<=signed(DIN_93_7)*signed(FMAP_32_93);
			MULT_94(31)<=signed(DIN_94_7)*signed(FMAP_32_94);
			MULT_95(31)<=signed(DIN_95_7)*signed(FMAP_32_95);
			MULT_96(31)<=signed(DIN_96_7)*signed(FMAP_32_96);
			MULT_97(31)<=signed(DIN_97_7)*signed(FMAP_32_97);
			MULT_98(31)<=signed(DIN_98_7)*signed(FMAP_32_98);
			MULT_99(31)<=signed(DIN_99_7)*signed(FMAP_32_99);
			MULT_100(31)<=signed(DIN_100_7)*signed(FMAP_32_100);
			MULT_101(31)<=signed(DIN_101_7)*signed(FMAP_32_101);
			MULT_102(31)<=signed(DIN_102_7)*signed(FMAP_32_102);
			MULT_103(31)<=signed(DIN_103_7)*signed(FMAP_32_103);
			MULT_104(31)<=signed(DIN_104_7)*signed(FMAP_32_104);
			MULT_105(31)<=signed(DIN_105_7)*signed(FMAP_32_105);
			MULT_106(31)<=signed(DIN_106_7)*signed(FMAP_32_106);
			MULT_107(31)<=signed(DIN_107_7)*signed(FMAP_32_107);
			MULT_108(31)<=signed(DIN_108_7)*signed(FMAP_32_108);
			MULT_109(31)<=signed(DIN_109_7)*signed(FMAP_32_109);
			MULT_110(31)<=signed(DIN_110_7)*signed(FMAP_32_110);
			MULT_111(31)<=signed(DIN_111_7)*signed(FMAP_32_111);
			MULT_112(31)<=signed(DIN_112_7)*signed(FMAP_32_112);
			MULT_113(31)<=signed(DIN_113_7)*signed(FMAP_32_113);
			MULT_114(31)<=signed(DIN_114_7)*signed(FMAP_32_114);
			MULT_115(31)<=signed(DIN_115_7)*signed(FMAP_32_115);
			MULT_116(31)<=signed(DIN_116_7)*signed(FMAP_32_116);
			MULT_117(31)<=signed(DIN_117_7)*signed(FMAP_32_117);
			MULT_118(31)<=signed(DIN_118_7)*signed(FMAP_32_118);
			MULT_119(31)<=signed(DIN_119_7)*signed(FMAP_32_119);
			MULT_120(31)<=signed(DIN_120_7)*signed(FMAP_32_120);

			MULT_1(32)<=signed(DIN_1_7)*signed(FMAP_33_1);
			MULT_2(32)<=signed(DIN_2_7)*signed(FMAP_33_2);
			MULT_3(32)<=signed(DIN_3_7)*signed(FMAP_33_3);
			MULT_4(32)<=signed(DIN_4_7)*signed(FMAP_33_4);
			MULT_5(32)<=signed(DIN_5_7)*signed(FMAP_33_5);
			MULT_6(32)<=signed(DIN_6_7)*signed(FMAP_33_6);
			MULT_7(32)<=signed(DIN_7_7)*signed(FMAP_33_7);
			MULT_8(32)<=signed(DIN_8_7)*signed(FMAP_33_8);
			MULT_9(32)<=signed(DIN_9_7)*signed(FMAP_33_9);
			MULT_10(32)<=signed(DIN_10_7)*signed(FMAP_33_10);
			MULT_11(32)<=signed(DIN_11_7)*signed(FMAP_33_11);
			MULT_12(32)<=signed(DIN_12_7)*signed(FMAP_33_12);
			MULT_13(32)<=signed(DIN_13_7)*signed(FMAP_33_13);
			MULT_14(32)<=signed(DIN_14_7)*signed(FMAP_33_14);
			MULT_15(32)<=signed(DIN_15_7)*signed(FMAP_33_15);
			MULT_16(32)<=signed(DIN_16_7)*signed(FMAP_33_16);
			MULT_17(32)<=signed(DIN_17_7)*signed(FMAP_33_17);
			MULT_18(32)<=signed(DIN_18_7)*signed(FMAP_33_18);
			MULT_19(32)<=signed(DIN_19_7)*signed(FMAP_33_19);
			MULT_20(32)<=signed(DIN_20_7)*signed(FMAP_33_20);
			MULT_21(32)<=signed(DIN_21_7)*signed(FMAP_33_21);
			MULT_22(32)<=signed(DIN_22_7)*signed(FMAP_33_22);
			MULT_23(32)<=signed(DIN_23_7)*signed(FMAP_33_23);
			MULT_24(32)<=signed(DIN_24_7)*signed(FMAP_33_24);
			MULT_25(32)<=signed(DIN_25_7)*signed(FMAP_33_25);
			MULT_26(32)<=signed(DIN_26_7)*signed(FMAP_33_26);
			MULT_27(32)<=signed(DIN_27_7)*signed(FMAP_33_27);
			MULT_28(32)<=signed(DIN_28_7)*signed(FMAP_33_28);
			MULT_29(32)<=signed(DIN_29_7)*signed(FMAP_33_29);
			MULT_30(32)<=signed(DIN_30_7)*signed(FMAP_33_30);
			MULT_31(32)<=signed(DIN_31_7)*signed(FMAP_33_31);
			MULT_32(32)<=signed(DIN_32_7)*signed(FMAP_33_32);
			MULT_33(32)<=signed(DIN_33_7)*signed(FMAP_33_33);
			MULT_34(32)<=signed(DIN_34_7)*signed(FMAP_33_34);
			MULT_35(32)<=signed(DIN_35_7)*signed(FMAP_33_35);
			MULT_36(32)<=signed(DIN_36_7)*signed(FMAP_33_36);
			MULT_37(32)<=signed(DIN_37_7)*signed(FMAP_33_37);
			MULT_38(32)<=signed(DIN_38_7)*signed(FMAP_33_38);
			MULT_39(32)<=signed(DIN_39_7)*signed(FMAP_33_39);
			MULT_40(32)<=signed(DIN_40_7)*signed(FMAP_33_40);
			MULT_41(32)<=signed(DIN_41_7)*signed(FMAP_33_41);
			MULT_42(32)<=signed(DIN_42_7)*signed(FMAP_33_42);
			MULT_43(32)<=signed(DIN_43_7)*signed(FMAP_33_43);
			MULT_44(32)<=signed(DIN_44_7)*signed(FMAP_33_44);
			MULT_45(32)<=signed(DIN_45_7)*signed(FMAP_33_45);
			MULT_46(32)<=signed(DIN_46_7)*signed(FMAP_33_46);
			MULT_47(32)<=signed(DIN_47_7)*signed(FMAP_33_47);
			MULT_48(32)<=signed(DIN_48_7)*signed(FMAP_33_48);
			MULT_49(32)<=signed(DIN_49_7)*signed(FMAP_33_49);
			MULT_50(32)<=signed(DIN_50_7)*signed(FMAP_33_50);
			MULT_51(32)<=signed(DIN_51_7)*signed(FMAP_33_51);
			MULT_52(32)<=signed(DIN_52_7)*signed(FMAP_33_52);
			MULT_53(32)<=signed(DIN_53_7)*signed(FMAP_33_53);
			MULT_54(32)<=signed(DIN_54_7)*signed(FMAP_33_54);
			MULT_55(32)<=signed(DIN_55_7)*signed(FMAP_33_55);
			MULT_56(32)<=signed(DIN_56_7)*signed(FMAP_33_56);
			MULT_57(32)<=signed(DIN_57_7)*signed(FMAP_33_57);
			MULT_58(32)<=signed(DIN_58_7)*signed(FMAP_33_58);
			MULT_59(32)<=signed(DIN_59_7)*signed(FMAP_33_59);
			MULT_60(32)<=signed(DIN_60_7)*signed(FMAP_33_60);
			MULT_61(32)<=signed(DIN_61_7)*signed(FMAP_33_61);
			MULT_62(32)<=signed(DIN_62_7)*signed(FMAP_33_62);
			MULT_63(32)<=signed(DIN_63_7)*signed(FMAP_33_63);
			MULT_64(32)<=signed(DIN_64_7)*signed(FMAP_33_64);
			MULT_65(32)<=signed(DIN_65_7)*signed(FMAP_33_65);
			MULT_66(32)<=signed(DIN_66_7)*signed(FMAP_33_66);
			MULT_67(32)<=signed(DIN_67_7)*signed(FMAP_33_67);
			MULT_68(32)<=signed(DIN_68_7)*signed(FMAP_33_68);
			MULT_69(32)<=signed(DIN_69_7)*signed(FMAP_33_69);
			MULT_70(32)<=signed(DIN_70_7)*signed(FMAP_33_70);
			MULT_71(32)<=signed(DIN_71_7)*signed(FMAP_33_71);
			MULT_72(32)<=signed(DIN_72_7)*signed(FMAP_33_72);
			MULT_73(32)<=signed(DIN_73_7)*signed(FMAP_33_73);
			MULT_74(32)<=signed(DIN_74_7)*signed(FMAP_33_74);
			MULT_75(32)<=signed(DIN_75_7)*signed(FMAP_33_75);
			MULT_76(32)<=signed(DIN_76_7)*signed(FMAP_33_76);
			MULT_77(32)<=signed(DIN_77_7)*signed(FMAP_33_77);
			MULT_78(32)<=signed(DIN_78_7)*signed(FMAP_33_78);
			MULT_79(32)<=signed(DIN_79_7)*signed(FMAP_33_79);
			MULT_80(32)<=signed(DIN_80_7)*signed(FMAP_33_80);
			MULT_81(32)<=signed(DIN_81_7)*signed(FMAP_33_81);
			MULT_82(32)<=signed(DIN_82_7)*signed(FMAP_33_82);
			MULT_83(32)<=signed(DIN_83_7)*signed(FMAP_33_83);
			MULT_84(32)<=signed(DIN_84_7)*signed(FMAP_33_84);
			MULT_85(32)<=signed(DIN_85_7)*signed(FMAP_33_85);
			MULT_86(32)<=signed(DIN_86_7)*signed(FMAP_33_86);
			MULT_87(32)<=signed(DIN_87_7)*signed(FMAP_33_87);
			MULT_88(32)<=signed(DIN_88_7)*signed(FMAP_33_88);
			MULT_89(32)<=signed(DIN_89_7)*signed(FMAP_33_89);
			MULT_90(32)<=signed(DIN_90_7)*signed(FMAP_33_90);
			MULT_91(32)<=signed(DIN_91_7)*signed(FMAP_33_91);
			MULT_92(32)<=signed(DIN_92_7)*signed(FMAP_33_92);
			MULT_93(32)<=signed(DIN_93_7)*signed(FMAP_33_93);
			MULT_94(32)<=signed(DIN_94_7)*signed(FMAP_33_94);
			MULT_95(32)<=signed(DIN_95_7)*signed(FMAP_33_95);
			MULT_96(32)<=signed(DIN_96_7)*signed(FMAP_33_96);
			MULT_97(32)<=signed(DIN_97_7)*signed(FMAP_33_97);
			MULT_98(32)<=signed(DIN_98_7)*signed(FMAP_33_98);
			MULT_99(32)<=signed(DIN_99_7)*signed(FMAP_33_99);
			MULT_100(32)<=signed(DIN_100_7)*signed(FMAP_33_100);
			MULT_101(32)<=signed(DIN_101_7)*signed(FMAP_33_101);
			MULT_102(32)<=signed(DIN_102_7)*signed(FMAP_33_102);
			MULT_103(32)<=signed(DIN_103_7)*signed(FMAP_33_103);
			MULT_104(32)<=signed(DIN_104_7)*signed(FMAP_33_104);
			MULT_105(32)<=signed(DIN_105_7)*signed(FMAP_33_105);
			MULT_106(32)<=signed(DIN_106_7)*signed(FMAP_33_106);
			MULT_107(32)<=signed(DIN_107_7)*signed(FMAP_33_107);
			MULT_108(32)<=signed(DIN_108_7)*signed(FMAP_33_108);
			MULT_109(32)<=signed(DIN_109_7)*signed(FMAP_33_109);
			MULT_110(32)<=signed(DIN_110_7)*signed(FMAP_33_110);
			MULT_111(32)<=signed(DIN_111_7)*signed(FMAP_33_111);
			MULT_112(32)<=signed(DIN_112_7)*signed(FMAP_33_112);
			MULT_113(32)<=signed(DIN_113_7)*signed(FMAP_33_113);
			MULT_114(32)<=signed(DIN_114_7)*signed(FMAP_33_114);
			MULT_115(32)<=signed(DIN_115_7)*signed(FMAP_33_115);
			MULT_116(32)<=signed(DIN_116_7)*signed(FMAP_33_116);
			MULT_117(32)<=signed(DIN_117_7)*signed(FMAP_33_117);
			MULT_118(32)<=signed(DIN_118_7)*signed(FMAP_33_118);
			MULT_119(32)<=signed(DIN_119_7)*signed(FMAP_33_119);
			MULT_120(32)<=signed(DIN_120_7)*signed(FMAP_33_120);

			MULT_1(33)<=signed(DIN_1_7)*signed(FMAP_34_1);
			MULT_2(33)<=signed(DIN_2_7)*signed(FMAP_34_2);
			MULT_3(33)<=signed(DIN_3_7)*signed(FMAP_34_3);
			MULT_4(33)<=signed(DIN_4_7)*signed(FMAP_34_4);
			MULT_5(33)<=signed(DIN_5_7)*signed(FMAP_34_5);
			MULT_6(33)<=signed(DIN_6_7)*signed(FMAP_34_6);
			MULT_7(33)<=signed(DIN_7_7)*signed(FMAP_34_7);
			MULT_8(33)<=signed(DIN_8_7)*signed(FMAP_34_8);
			MULT_9(33)<=signed(DIN_9_7)*signed(FMAP_34_9);
			MULT_10(33)<=signed(DIN_10_7)*signed(FMAP_34_10);
			MULT_11(33)<=signed(DIN_11_7)*signed(FMAP_34_11);
			MULT_12(33)<=signed(DIN_12_7)*signed(FMAP_34_12);
			MULT_13(33)<=signed(DIN_13_7)*signed(FMAP_34_13);
			MULT_14(33)<=signed(DIN_14_7)*signed(FMAP_34_14);
			MULT_15(33)<=signed(DIN_15_7)*signed(FMAP_34_15);
			MULT_16(33)<=signed(DIN_16_7)*signed(FMAP_34_16);
			MULT_17(33)<=signed(DIN_17_7)*signed(FMAP_34_17);
			MULT_18(33)<=signed(DIN_18_7)*signed(FMAP_34_18);
			MULT_19(33)<=signed(DIN_19_7)*signed(FMAP_34_19);
			MULT_20(33)<=signed(DIN_20_7)*signed(FMAP_34_20);
			MULT_21(33)<=signed(DIN_21_7)*signed(FMAP_34_21);
			MULT_22(33)<=signed(DIN_22_7)*signed(FMAP_34_22);
			MULT_23(33)<=signed(DIN_23_7)*signed(FMAP_34_23);
			MULT_24(33)<=signed(DIN_24_7)*signed(FMAP_34_24);
			MULT_25(33)<=signed(DIN_25_7)*signed(FMAP_34_25);
			MULT_26(33)<=signed(DIN_26_7)*signed(FMAP_34_26);
			MULT_27(33)<=signed(DIN_27_7)*signed(FMAP_34_27);
			MULT_28(33)<=signed(DIN_28_7)*signed(FMAP_34_28);
			MULT_29(33)<=signed(DIN_29_7)*signed(FMAP_34_29);
			MULT_30(33)<=signed(DIN_30_7)*signed(FMAP_34_30);
			MULT_31(33)<=signed(DIN_31_7)*signed(FMAP_34_31);
			MULT_32(33)<=signed(DIN_32_7)*signed(FMAP_34_32);
			MULT_33(33)<=signed(DIN_33_7)*signed(FMAP_34_33);
			MULT_34(33)<=signed(DIN_34_7)*signed(FMAP_34_34);
			MULT_35(33)<=signed(DIN_35_7)*signed(FMAP_34_35);
			MULT_36(33)<=signed(DIN_36_7)*signed(FMAP_34_36);
			MULT_37(33)<=signed(DIN_37_7)*signed(FMAP_34_37);
			MULT_38(33)<=signed(DIN_38_7)*signed(FMAP_34_38);
			MULT_39(33)<=signed(DIN_39_7)*signed(FMAP_34_39);
			MULT_40(33)<=signed(DIN_40_7)*signed(FMAP_34_40);
			MULT_41(33)<=signed(DIN_41_7)*signed(FMAP_34_41);
			MULT_42(33)<=signed(DIN_42_7)*signed(FMAP_34_42);
			MULT_43(33)<=signed(DIN_43_7)*signed(FMAP_34_43);
			MULT_44(33)<=signed(DIN_44_7)*signed(FMAP_34_44);
			MULT_45(33)<=signed(DIN_45_7)*signed(FMAP_34_45);
			MULT_46(33)<=signed(DIN_46_7)*signed(FMAP_34_46);
			MULT_47(33)<=signed(DIN_47_7)*signed(FMAP_34_47);
			MULT_48(33)<=signed(DIN_48_7)*signed(FMAP_34_48);
			MULT_49(33)<=signed(DIN_49_7)*signed(FMAP_34_49);
			MULT_50(33)<=signed(DIN_50_7)*signed(FMAP_34_50);
			MULT_51(33)<=signed(DIN_51_7)*signed(FMAP_34_51);
			MULT_52(33)<=signed(DIN_52_7)*signed(FMAP_34_52);
			MULT_53(33)<=signed(DIN_53_7)*signed(FMAP_34_53);
			MULT_54(33)<=signed(DIN_54_7)*signed(FMAP_34_54);
			MULT_55(33)<=signed(DIN_55_7)*signed(FMAP_34_55);
			MULT_56(33)<=signed(DIN_56_7)*signed(FMAP_34_56);
			MULT_57(33)<=signed(DIN_57_7)*signed(FMAP_34_57);
			MULT_58(33)<=signed(DIN_58_7)*signed(FMAP_34_58);
			MULT_59(33)<=signed(DIN_59_7)*signed(FMAP_34_59);
			MULT_60(33)<=signed(DIN_60_7)*signed(FMAP_34_60);
			MULT_61(33)<=signed(DIN_61_7)*signed(FMAP_34_61);
			MULT_62(33)<=signed(DIN_62_7)*signed(FMAP_34_62);
			MULT_63(33)<=signed(DIN_63_7)*signed(FMAP_34_63);
			MULT_64(33)<=signed(DIN_64_7)*signed(FMAP_34_64);
			MULT_65(33)<=signed(DIN_65_7)*signed(FMAP_34_65);
			MULT_66(33)<=signed(DIN_66_7)*signed(FMAP_34_66);
			MULT_67(33)<=signed(DIN_67_7)*signed(FMAP_34_67);
			MULT_68(33)<=signed(DIN_68_7)*signed(FMAP_34_68);
			MULT_69(33)<=signed(DIN_69_7)*signed(FMAP_34_69);
			MULT_70(33)<=signed(DIN_70_7)*signed(FMAP_34_70);
			MULT_71(33)<=signed(DIN_71_7)*signed(FMAP_34_71);
			MULT_72(33)<=signed(DIN_72_7)*signed(FMAP_34_72);
			MULT_73(33)<=signed(DIN_73_7)*signed(FMAP_34_73);
			MULT_74(33)<=signed(DIN_74_7)*signed(FMAP_34_74);
			MULT_75(33)<=signed(DIN_75_7)*signed(FMAP_34_75);
			MULT_76(33)<=signed(DIN_76_7)*signed(FMAP_34_76);
			MULT_77(33)<=signed(DIN_77_7)*signed(FMAP_34_77);
			MULT_78(33)<=signed(DIN_78_7)*signed(FMAP_34_78);
			MULT_79(33)<=signed(DIN_79_7)*signed(FMAP_34_79);
			MULT_80(33)<=signed(DIN_80_7)*signed(FMAP_34_80);
			MULT_81(33)<=signed(DIN_81_7)*signed(FMAP_34_81);
			MULT_82(33)<=signed(DIN_82_7)*signed(FMAP_34_82);
			MULT_83(33)<=signed(DIN_83_7)*signed(FMAP_34_83);
			MULT_84(33)<=signed(DIN_84_7)*signed(FMAP_34_84);
			MULT_85(33)<=signed(DIN_85_7)*signed(FMAP_34_85);
			MULT_86(33)<=signed(DIN_86_7)*signed(FMAP_34_86);
			MULT_87(33)<=signed(DIN_87_7)*signed(FMAP_34_87);
			MULT_88(33)<=signed(DIN_88_7)*signed(FMAP_34_88);
			MULT_89(33)<=signed(DIN_89_7)*signed(FMAP_34_89);
			MULT_90(33)<=signed(DIN_90_7)*signed(FMAP_34_90);
			MULT_91(33)<=signed(DIN_91_7)*signed(FMAP_34_91);
			MULT_92(33)<=signed(DIN_92_7)*signed(FMAP_34_92);
			MULT_93(33)<=signed(DIN_93_7)*signed(FMAP_34_93);
			MULT_94(33)<=signed(DIN_94_7)*signed(FMAP_34_94);
			MULT_95(33)<=signed(DIN_95_7)*signed(FMAP_34_95);
			MULT_96(33)<=signed(DIN_96_7)*signed(FMAP_34_96);
			MULT_97(33)<=signed(DIN_97_7)*signed(FMAP_34_97);
			MULT_98(33)<=signed(DIN_98_7)*signed(FMAP_34_98);
			MULT_99(33)<=signed(DIN_99_7)*signed(FMAP_34_99);
			MULT_100(33)<=signed(DIN_100_7)*signed(FMAP_34_100);
			MULT_101(33)<=signed(DIN_101_7)*signed(FMAP_34_101);
			MULT_102(33)<=signed(DIN_102_7)*signed(FMAP_34_102);
			MULT_103(33)<=signed(DIN_103_7)*signed(FMAP_34_103);
			MULT_104(33)<=signed(DIN_104_7)*signed(FMAP_34_104);
			MULT_105(33)<=signed(DIN_105_7)*signed(FMAP_34_105);
			MULT_106(33)<=signed(DIN_106_7)*signed(FMAP_34_106);
			MULT_107(33)<=signed(DIN_107_7)*signed(FMAP_34_107);
			MULT_108(33)<=signed(DIN_108_7)*signed(FMAP_34_108);
			MULT_109(33)<=signed(DIN_109_7)*signed(FMAP_34_109);
			MULT_110(33)<=signed(DIN_110_7)*signed(FMAP_34_110);
			MULT_111(33)<=signed(DIN_111_7)*signed(FMAP_34_111);
			MULT_112(33)<=signed(DIN_112_7)*signed(FMAP_34_112);
			MULT_113(33)<=signed(DIN_113_7)*signed(FMAP_34_113);
			MULT_114(33)<=signed(DIN_114_7)*signed(FMAP_34_114);
			MULT_115(33)<=signed(DIN_115_7)*signed(FMAP_34_115);
			MULT_116(33)<=signed(DIN_116_7)*signed(FMAP_34_116);
			MULT_117(33)<=signed(DIN_117_7)*signed(FMAP_34_117);
			MULT_118(33)<=signed(DIN_118_7)*signed(FMAP_34_118);
			MULT_119(33)<=signed(DIN_119_7)*signed(FMAP_34_119);
			MULT_120(33)<=signed(DIN_120_7)*signed(FMAP_34_120);

			MULT_1(34)<=signed(DIN_1_7)*signed(FMAP_35_1);
			MULT_2(34)<=signed(DIN_2_7)*signed(FMAP_35_2);
			MULT_3(34)<=signed(DIN_3_7)*signed(FMAP_35_3);
			MULT_4(34)<=signed(DIN_4_7)*signed(FMAP_35_4);
			MULT_5(34)<=signed(DIN_5_7)*signed(FMAP_35_5);
			MULT_6(34)<=signed(DIN_6_7)*signed(FMAP_35_6);
			MULT_7(34)<=signed(DIN_7_7)*signed(FMAP_35_7);
			MULT_8(34)<=signed(DIN_8_7)*signed(FMAP_35_8);
			MULT_9(34)<=signed(DIN_9_7)*signed(FMAP_35_9);
			MULT_10(34)<=signed(DIN_10_7)*signed(FMAP_35_10);
			MULT_11(34)<=signed(DIN_11_7)*signed(FMAP_35_11);
			MULT_12(34)<=signed(DIN_12_7)*signed(FMAP_35_12);
			MULT_13(34)<=signed(DIN_13_7)*signed(FMAP_35_13);
			MULT_14(34)<=signed(DIN_14_7)*signed(FMAP_35_14);
			MULT_15(34)<=signed(DIN_15_7)*signed(FMAP_35_15);
			MULT_16(34)<=signed(DIN_16_7)*signed(FMAP_35_16);
			MULT_17(34)<=signed(DIN_17_7)*signed(FMAP_35_17);
			MULT_18(34)<=signed(DIN_18_7)*signed(FMAP_35_18);
			MULT_19(34)<=signed(DIN_19_7)*signed(FMAP_35_19);
			MULT_20(34)<=signed(DIN_20_7)*signed(FMAP_35_20);
			MULT_21(34)<=signed(DIN_21_7)*signed(FMAP_35_21);
			MULT_22(34)<=signed(DIN_22_7)*signed(FMAP_35_22);
			MULT_23(34)<=signed(DIN_23_7)*signed(FMAP_35_23);
			MULT_24(34)<=signed(DIN_24_7)*signed(FMAP_35_24);
			MULT_25(34)<=signed(DIN_25_7)*signed(FMAP_35_25);
			MULT_26(34)<=signed(DIN_26_7)*signed(FMAP_35_26);
			MULT_27(34)<=signed(DIN_27_7)*signed(FMAP_35_27);
			MULT_28(34)<=signed(DIN_28_7)*signed(FMAP_35_28);
			MULT_29(34)<=signed(DIN_29_7)*signed(FMAP_35_29);
			MULT_30(34)<=signed(DIN_30_7)*signed(FMAP_35_30);
			MULT_31(34)<=signed(DIN_31_7)*signed(FMAP_35_31);
			MULT_32(34)<=signed(DIN_32_7)*signed(FMAP_35_32);
			MULT_33(34)<=signed(DIN_33_7)*signed(FMAP_35_33);
			MULT_34(34)<=signed(DIN_34_7)*signed(FMAP_35_34);
			MULT_35(34)<=signed(DIN_35_7)*signed(FMAP_35_35);
			MULT_36(34)<=signed(DIN_36_7)*signed(FMAP_35_36);
			MULT_37(34)<=signed(DIN_37_7)*signed(FMAP_35_37);
			MULT_38(34)<=signed(DIN_38_7)*signed(FMAP_35_38);
			MULT_39(34)<=signed(DIN_39_7)*signed(FMAP_35_39);
			MULT_40(34)<=signed(DIN_40_7)*signed(FMAP_35_40);
			MULT_41(34)<=signed(DIN_41_7)*signed(FMAP_35_41);
			MULT_42(34)<=signed(DIN_42_7)*signed(FMAP_35_42);
			MULT_43(34)<=signed(DIN_43_7)*signed(FMAP_35_43);
			MULT_44(34)<=signed(DIN_44_7)*signed(FMAP_35_44);
			MULT_45(34)<=signed(DIN_45_7)*signed(FMAP_35_45);
			MULT_46(34)<=signed(DIN_46_7)*signed(FMAP_35_46);
			MULT_47(34)<=signed(DIN_47_7)*signed(FMAP_35_47);
			MULT_48(34)<=signed(DIN_48_7)*signed(FMAP_35_48);
			MULT_49(34)<=signed(DIN_49_7)*signed(FMAP_35_49);
			MULT_50(34)<=signed(DIN_50_7)*signed(FMAP_35_50);
			MULT_51(34)<=signed(DIN_51_7)*signed(FMAP_35_51);
			MULT_52(34)<=signed(DIN_52_7)*signed(FMAP_35_52);
			MULT_53(34)<=signed(DIN_53_7)*signed(FMAP_35_53);
			MULT_54(34)<=signed(DIN_54_7)*signed(FMAP_35_54);
			MULT_55(34)<=signed(DIN_55_7)*signed(FMAP_35_55);
			MULT_56(34)<=signed(DIN_56_7)*signed(FMAP_35_56);
			MULT_57(34)<=signed(DIN_57_7)*signed(FMAP_35_57);
			MULT_58(34)<=signed(DIN_58_7)*signed(FMAP_35_58);
			MULT_59(34)<=signed(DIN_59_7)*signed(FMAP_35_59);
			MULT_60(34)<=signed(DIN_60_7)*signed(FMAP_35_60);
			MULT_61(34)<=signed(DIN_61_7)*signed(FMAP_35_61);
			MULT_62(34)<=signed(DIN_62_7)*signed(FMAP_35_62);
			MULT_63(34)<=signed(DIN_63_7)*signed(FMAP_35_63);
			MULT_64(34)<=signed(DIN_64_7)*signed(FMAP_35_64);
			MULT_65(34)<=signed(DIN_65_7)*signed(FMAP_35_65);
			MULT_66(34)<=signed(DIN_66_7)*signed(FMAP_35_66);
			MULT_67(34)<=signed(DIN_67_7)*signed(FMAP_35_67);
			MULT_68(34)<=signed(DIN_68_7)*signed(FMAP_35_68);
			MULT_69(34)<=signed(DIN_69_7)*signed(FMAP_35_69);
			MULT_70(34)<=signed(DIN_70_7)*signed(FMAP_35_70);
			MULT_71(34)<=signed(DIN_71_7)*signed(FMAP_35_71);
			MULT_72(34)<=signed(DIN_72_7)*signed(FMAP_35_72);
			MULT_73(34)<=signed(DIN_73_7)*signed(FMAP_35_73);
			MULT_74(34)<=signed(DIN_74_7)*signed(FMAP_35_74);
			MULT_75(34)<=signed(DIN_75_7)*signed(FMAP_35_75);
			MULT_76(34)<=signed(DIN_76_7)*signed(FMAP_35_76);
			MULT_77(34)<=signed(DIN_77_7)*signed(FMAP_35_77);
			MULT_78(34)<=signed(DIN_78_7)*signed(FMAP_35_78);
			MULT_79(34)<=signed(DIN_79_7)*signed(FMAP_35_79);
			MULT_80(34)<=signed(DIN_80_7)*signed(FMAP_35_80);
			MULT_81(34)<=signed(DIN_81_7)*signed(FMAP_35_81);
			MULT_82(34)<=signed(DIN_82_7)*signed(FMAP_35_82);
			MULT_83(34)<=signed(DIN_83_7)*signed(FMAP_35_83);
			MULT_84(34)<=signed(DIN_84_7)*signed(FMAP_35_84);
			MULT_85(34)<=signed(DIN_85_7)*signed(FMAP_35_85);
			MULT_86(34)<=signed(DIN_86_7)*signed(FMAP_35_86);
			MULT_87(34)<=signed(DIN_87_7)*signed(FMAP_35_87);
			MULT_88(34)<=signed(DIN_88_7)*signed(FMAP_35_88);
			MULT_89(34)<=signed(DIN_89_7)*signed(FMAP_35_89);
			MULT_90(34)<=signed(DIN_90_7)*signed(FMAP_35_90);
			MULT_91(34)<=signed(DIN_91_7)*signed(FMAP_35_91);
			MULT_92(34)<=signed(DIN_92_7)*signed(FMAP_35_92);
			MULT_93(34)<=signed(DIN_93_7)*signed(FMAP_35_93);
			MULT_94(34)<=signed(DIN_94_7)*signed(FMAP_35_94);
			MULT_95(34)<=signed(DIN_95_7)*signed(FMAP_35_95);
			MULT_96(34)<=signed(DIN_96_7)*signed(FMAP_35_96);
			MULT_97(34)<=signed(DIN_97_7)*signed(FMAP_35_97);
			MULT_98(34)<=signed(DIN_98_7)*signed(FMAP_35_98);
			MULT_99(34)<=signed(DIN_99_7)*signed(FMAP_35_99);
			MULT_100(34)<=signed(DIN_100_7)*signed(FMAP_35_100);
			MULT_101(34)<=signed(DIN_101_7)*signed(FMAP_35_101);
			MULT_102(34)<=signed(DIN_102_7)*signed(FMAP_35_102);
			MULT_103(34)<=signed(DIN_103_7)*signed(FMAP_35_103);
			MULT_104(34)<=signed(DIN_104_7)*signed(FMAP_35_104);
			MULT_105(34)<=signed(DIN_105_7)*signed(FMAP_35_105);
			MULT_106(34)<=signed(DIN_106_7)*signed(FMAP_35_106);
			MULT_107(34)<=signed(DIN_107_7)*signed(FMAP_35_107);
			MULT_108(34)<=signed(DIN_108_7)*signed(FMAP_35_108);
			MULT_109(34)<=signed(DIN_109_7)*signed(FMAP_35_109);
			MULT_110(34)<=signed(DIN_110_7)*signed(FMAP_35_110);
			MULT_111(34)<=signed(DIN_111_7)*signed(FMAP_35_111);
			MULT_112(34)<=signed(DIN_112_7)*signed(FMAP_35_112);
			MULT_113(34)<=signed(DIN_113_7)*signed(FMAP_35_113);
			MULT_114(34)<=signed(DIN_114_7)*signed(FMAP_35_114);
			MULT_115(34)<=signed(DIN_115_7)*signed(FMAP_35_115);
			MULT_116(34)<=signed(DIN_116_7)*signed(FMAP_35_116);
			MULT_117(34)<=signed(DIN_117_7)*signed(FMAP_35_117);
			MULT_118(34)<=signed(DIN_118_7)*signed(FMAP_35_118);
			MULT_119(34)<=signed(DIN_119_7)*signed(FMAP_35_119);
			MULT_120(34)<=signed(DIN_120_7)*signed(FMAP_35_120);

			MULT_1(35)<=signed(DIN_1_7)*signed(FMAP_36_1);
			MULT_2(35)<=signed(DIN_2_7)*signed(FMAP_36_2);
			MULT_3(35)<=signed(DIN_3_7)*signed(FMAP_36_3);
			MULT_4(35)<=signed(DIN_4_7)*signed(FMAP_36_4);
			MULT_5(35)<=signed(DIN_5_7)*signed(FMAP_36_5);
			MULT_6(35)<=signed(DIN_6_7)*signed(FMAP_36_6);
			MULT_7(35)<=signed(DIN_7_7)*signed(FMAP_36_7);
			MULT_8(35)<=signed(DIN_8_7)*signed(FMAP_36_8);
			MULT_9(35)<=signed(DIN_9_7)*signed(FMAP_36_9);
			MULT_10(35)<=signed(DIN_10_7)*signed(FMAP_36_10);
			MULT_11(35)<=signed(DIN_11_7)*signed(FMAP_36_11);
			MULT_12(35)<=signed(DIN_12_7)*signed(FMAP_36_12);
			MULT_13(35)<=signed(DIN_13_7)*signed(FMAP_36_13);
			MULT_14(35)<=signed(DIN_14_7)*signed(FMAP_36_14);
			MULT_15(35)<=signed(DIN_15_7)*signed(FMAP_36_15);
			MULT_16(35)<=signed(DIN_16_7)*signed(FMAP_36_16);
			MULT_17(35)<=signed(DIN_17_7)*signed(FMAP_36_17);
			MULT_18(35)<=signed(DIN_18_7)*signed(FMAP_36_18);
			MULT_19(35)<=signed(DIN_19_7)*signed(FMAP_36_19);
			MULT_20(35)<=signed(DIN_20_7)*signed(FMAP_36_20);
			MULT_21(35)<=signed(DIN_21_7)*signed(FMAP_36_21);
			MULT_22(35)<=signed(DIN_22_7)*signed(FMAP_36_22);
			MULT_23(35)<=signed(DIN_23_7)*signed(FMAP_36_23);
			MULT_24(35)<=signed(DIN_24_7)*signed(FMAP_36_24);
			MULT_25(35)<=signed(DIN_25_7)*signed(FMAP_36_25);
			MULT_26(35)<=signed(DIN_26_7)*signed(FMAP_36_26);
			MULT_27(35)<=signed(DIN_27_7)*signed(FMAP_36_27);
			MULT_28(35)<=signed(DIN_28_7)*signed(FMAP_36_28);
			MULT_29(35)<=signed(DIN_29_7)*signed(FMAP_36_29);
			MULT_30(35)<=signed(DIN_30_7)*signed(FMAP_36_30);
			MULT_31(35)<=signed(DIN_31_7)*signed(FMAP_36_31);
			MULT_32(35)<=signed(DIN_32_7)*signed(FMAP_36_32);
			MULT_33(35)<=signed(DIN_33_7)*signed(FMAP_36_33);
			MULT_34(35)<=signed(DIN_34_7)*signed(FMAP_36_34);
			MULT_35(35)<=signed(DIN_35_7)*signed(FMAP_36_35);
			MULT_36(35)<=signed(DIN_36_7)*signed(FMAP_36_36);
			MULT_37(35)<=signed(DIN_37_7)*signed(FMAP_36_37);
			MULT_38(35)<=signed(DIN_38_7)*signed(FMAP_36_38);
			MULT_39(35)<=signed(DIN_39_7)*signed(FMAP_36_39);
			MULT_40(35)<=signed(DIN_40_7)*signed(FMAP_36_40);
			MULT_41(35)<=signed(DIN_41_7)*signed(FMAP_36_41);
			MULT_42(35)<=signed(DIN_42_7)*signed(FMAP_36_42);
			MULT_43(35)<=signed(DIN_43_7)*signed(FMAP_36_43);
			MULT_44(35)<=signed(DIN_44_7)*signed(FMAP_36_44);
			MULT_45(35)<=signed(DIN_45_7)*signed(FMAP_36_45);
			MULT_46(35)<=signed(DIN_46_7)*signed(FMAP_36_46);
			MULT_47(35)<=signed(DIN_47_7)*signed(FMAP_36_47);
			MULT_48(35)<=signed(DIN_48_7)*signed(FMAP_36_48);
			MULT_49(35)<=signed(DIN_49_7)*signed(FMAP_36_49);
			MULT_50(35)<=signed(DIN_50_7)*signed(FMAP_36_50);
			MULT_51(35)<=signed(DIN_51_7)*signed(FMAP_36_51);
			MULT_52(35)<=signed(DIN_52_7)*signed(FMAP_36_52);
			MULT_53(35)<=signed(DIN_53_7)*signed(FMAP_36_53);
			MULT_54(35)<=signed(DIN_54_7)*signed(FMAP_36_54);
			MULT_55(35)<=signed(DIN_55_7)*signed(FMAP_36_55);
			MULT_56(35)<=signed(DIN_56_7)*signed(FMAP_36_56);
			MULT_57(35)<=signed(DIN_57_7)*signed(FMAP_36_57);
			MULT_58(35)<=signed(DIN_58_7)*signed(FMAP_36_58);
			MULT_59(35)<=signed(DIN_59_7)*signed(FMAP_36_59);
			MULT_60(35)<=signed(DIN_60_7)*signed(FMAP_36_60);
			MULT_61(35)<=signed(DIN_61_7)*signed(FMAP_36_61);
			MULT_62(35)<=signed(DIN_62_7)*signed(FMAP_36_62);
			MULT_63(35)<=signed(DIN_63_7)*signed(FMAP_36_63);
			MULT_64(35)<=signed(DIN_64_7)*signed(FMAP_36_64);
			MULT_65(35)<=signed(DIN_65_7)*signed(FMAP_36_65);
			MULT_66(35)<=signed(DIN_66_7)*signed(FMAP_36_66);
			MULT_67(35)<=signed(DIN_67_7)*signed(FMAP_36_67);
			MULT_68(35)<=signed(DIN_68_7)*signed(FMAP_36_68);
			MULT_69(35)<=signed(DIN_69_7)*signed(FMAP_36_69);
			MULT_70(35)<=signed(DIN_70_7)*signed(FMAP_36_70);
			MULT_71(35)<=signed(DIN_71_7)*signed(FMAP_36_71);
			MULT_72(35)<=signed(DIN_72_7)*signed(FMAP_36_72);
			MULT_73(35)<=signed(DIN_73_7)*signed(FMAP_36_73);
			MULT_74(35)<=signed(DIN_74_7)*signed(FMAP_36_74);
			MULT_75(35)<=signed(DIN_75_7)*signed(FMAP_36_75);
			MULT_76(35)<=signed(DIN_76_7)*signed(FMAP_36_76);
			MULT_77(35)<=signed(DIN_77_7)*signed(FMAP_36_77);
			MULT_78(35)<=signed(DIN_78_7)*signed(FMAP_36_78);
			MULT_79(35)<=signed(DIN_79_7)*signed(FMAP_36_79);
			MULT_80(35)<=signed(DIN_80_7)*signed(FMAP_36_80);
			MULT_81(35)<=signed(DIN_81_7)*signed(FMAP_36_81);
			MULT_82(35)<=signed(DIN_82_7)*signed(FMAP_36_82);
			MULT_83(35)<=signed(DIN_83_7)*signed(FMAP_36_83);
			MULT_84(35)<=signed(DIN_84_7)*signed(FMAP_36_84);
			MULT_85(35)<=signed(DIN_85_7)*signed(FMAP_36_85);
			MULT_86(35)<=signed(DIN_86_7)*signed(FMAP_36_86);
			MULT_87(35)<=signed(DIN_87_7)*signed(FMAP_36_87);
			MULT_88(35)<=signed(DIN_88_7)*signed(FMAP_36_88);
			MULT_89(35)<=signed(DIN_89_7)*signed(FMAP_36_89);
			MULT_90(35)<=signed(DIN_90_7)*signed(FMAP_36_90);
			MULT_91(35)<=signed(DIN_91_7)*signed(FMAP_36_91);
			MULT_92(35)<=signed(DIN_92_7)*signed(FMAP_36_92);
			MULT_93(35)<=signed(DIN_93_7)*signed(FMAP_36_93);
			MULT_94(35)<=signed(DIN_94_7)*signed(FMAP_36_94);
			MULT_95(35)<=signed(DIN_95_7)*signed(FMAP_36_95);
			MULT_96(35)<=signed(DIN_96_7)*signed(FMAP_36_96);
			MULT_97(35)<=signed(DIN_97_7)*signed(FMAP_36_97);
			MULT_98(35)<=signed(DIN_98_7)*signed(FMAP_36_98);
			MULT_99(35)<=signed(DIN_99_7)*signed(FMAP_36_99);
			MULT_100(35)<=signed(DIN_100_7)*signed(FMAP_36_100);
			MULT_101(35)<=signed(DIN_101_7)*signed(FMAP_36_101);
			MULT_102(35)<=signed(DIN_102_7)*signed(FMAP_36_102);
			MULT_103(35)<=signed(DIN_103_7)*signed(FMAP_36_103);
			MULT_104(35)<=signed(DIN_104_7)*signed(FMAP_36_104);
			MULT_105(35)<=signed(DIN_105_7)*signed(FMAP_36_105);
			MULT_106(35)<=signed(DIN_106_7)*signed(FMAP_36_106);
			MULT_107(35)<=signed(DIN_107_7)*signed(FMAP_36_107);
			MULT_108(35)<=signed(DIN_108_7)*signed(FMAP_36_108);
			MULT_109(35)<=signed(DIN_109_7)*signed(FMAP_36_109);
			MULT_110(35)<=signed(DIN_110_7)*signed(FMAP_36_110);
			MULT_111(35)<=signed(DIN_111_7)*signed(FMAP_36_111);
			MULT_112(35)<=signed(DIN_112_7)*signed(FMAP_36_112);
			MULT_113(35)<=signed(DIN_113_7)*signed(FMAP_36_113);
			MULT_114(35)<=signed(DIN_114_7)*signed(FMAP_36_114);
			MULT_115(35)<=signed(DIN_115_7)*signed(FMAP_36_115);
			MULT_116(35)<=signed(DIN_116_7)*signed(FMAP_36_116);
			MULT_117(35)<=signed(DIN_117_7)*signed(FMAP_36_117);
			MULT_118(35)<=signed(DIN_118_7)*signed(FMAP_36_118);
			MULT_119(35)<=signed(DIN_119_7)*signed(FMAP_36_119);
			MULT_120(35)<=signed(DIN_120_7)*signed(FMAP_36_120);

			MULT_1(36)<=signed(DIN_1_7)*signed(FMAP_37_1);
			MULT_2(36)<=signed(DIN_2_7)*signed(FMAP_37_2);
			MULT_3(36)<=signed(DIN_3_7)*signed(FMAP_37_3);
			MULT_4(36)<=signed(DIN_4_7)*signed(FMAP_37_4);
			MULT_5(36)<=signed(DIN_5_7)*signed(FMAP_37_5);
			MULT_6(36)<=signed(DIN_6_7)*signed(FMAP_37_6);
			MULT_7(36)<=signed(DIN_7_7)*signed(FMAP_37_7);
			MULT_8(36)<=signed(DIN_8_7)*signed(FMAP_37_8);
			MULT_9(36)<=signed(DIN_9_7)*signed(FMAP_37_9);
			MULT_10(36)<=signed(DIN_10_7)*signed(FMAP_37_10);
			MULT_11(36)<=signed(DIN_11_7)*signed(FMAP_37_11);
			MULT_12(36)<=signed(DIN_12_7)*signed(FMAP_37_12);
			MULT_13(36)<=signed(DIN_13_7)*signed(FMAP_37_13);
			MULT_14(36)<=signed(DIN_14_7)*signed(FMAP_37_14);
			MULT_15(36)<=signed(DIN_15_7)*signed(FMAP_37_15);
			MULT_16(36)<=signed(DIN_16_7)*signed(FMAP_37_16);
			MULT_17(36)<=signed(DIN_17_7)*signed(FMAP_37_17);
			MULT_18(36)<=signed(DIN_18_7)*signed(FMAP_37_18);
			MULT_19(36)<=signed(DIN_19_7)*signed(FMAP_37_19);
			MULT_20(36)<=signed(DIN_20_7)*signed(FMAP_37_20);
			MULT_21(36)<=signed(DIN_21_7)*signed(FMAP_37_21);
			MULT_22(36)<=signed(DIN_22_7)*signed(FMAP_37_22);
			MULT_23(36)<=signed(DIN_23_7)*signed(FMAP_37_23);
			MULT_24(36)<=signed(DIN_24_7)*signed(FMAP_37_24);
			MULT_25(36)<=signed(DIN_25_7)*signed(FMAP_37_25);
			MULT_26(36)<=signed(DIN_26_7)*signed(FMAP_37_26);
			MULT_27(36)<=signed(DIN_27_7)*signed(FMAP_37_27);
			MULT_28(36)<=signed(DIN_28_7)*signed(FMAP_37_28);
			MULT_29(36)<=signed(DIN_29_7)*signed(FMAP_37_29);
			MULT_30(36)<=signed(DIN_30_7)*signed(FMAP_37_30);
			MULT_31(36)<=signed(DIN_31_7)*signed(FMAP_37_31);
			MULT_32(36)<=signed(DIN_32_7)*signed(FMAP_37_32);
			MULT_33(36)<=signed(DIN_33_7)*signed(FMAP_37_33);
			MULT_34(36)<=signed(DIN_34_7)*signed(FMAP_37_34);
			MULT_35(36)<=signed(DIN_35_7)*signed(FMAP_37_35);
			MULT_36(36)<=signed(DIN_36_7)*signed(FMAP_37_36);
			MULT_37(36)<=signed(DIN_37_7)*signed(FMAP_37_37);
			MULT_38(36)<=signed(DIN_38_7)*signed(FMAP_37_38);
			MULT_39(36)<=signed(DIN_39_7)*signed(FMAP_37_39);
			MULT_40(36)<=signed(DIN_40_7)*signed(FMAP_37_40);
			MULT_41(36)<=signed(DIN_41_7)*signed(FMAP_37_41);
			MULT_42(36)<=signed(DIN_42_7)*signed(FMAP_37_42);
			MULT_43(36)<=signed(DIN_43_7)*signed(FMAP_37_43);
			MULT_44(36)<=signed(DIN_44_7)*signed(FMAP_37_44);
			MULT_45(36)<=signed(DIN_45_7)*signed(FMAP_37_45);
			MULT_46(36)<=signed(DIN_46_7)*signed(FMAP_37_46);
			MULT_47(36)<=signed(DIN_47_7)*signed(FMAP_37_47);
			MULT_48(36)<=signed(DIN_48_7)*signed(FMAP_37_48);
			MULT_49(36)<=signed(DIN_49_7)*signed(FMAP_37_49);
			MULT_50(36)<=signed(DIN_50_7)*signed(FMAP_37_50);
			MULT_51(36)<=signed(DIN_51_7)*signed(FMAP_37_51);
			MULT_52(36)<=signed(DIN_52_7)*signed(FMAP_37_52);
			MULT_53(36)<=signed(DIN_53_7)*signed(FMAP_37_53);
			MULT_54(36)<=signed(DIN_54_7)*signed(FMAP_37_54);
			MULT_55(36)<=signed(DIN_55_7)*signed(FMAP_37_55);
			MULT_56(36)<=signed(DIN_56_7)*signed(FMAP_37_56);
			MULT_57(36)<=signed(DIN_57_7)*signed(FMAP_37_57);
			MULT_58(36)<=signed(DIN_58_7)*signed(FMAP_37_58);
			MULT_59(36)<=signed(DIN_59_7)*signed(FMAP_37_59);
			MULT_60(36)<=signed(DIN_60_7)*signed(FMAP_37_60);
			MULT_61(36)<=signed(DIN_61_7)*signed(FMAP_37_61);
			MULT_62(36)<=signed(DIN_62_7)*signed(FMAP_37_62);
			MULT_63(36)<=signed(DIN_63_7)*signed(FMAP_37_63);
			MULT_64(36)<=signed(DIN_64_7)*signed(FMAP_37_64);
			MULT_65(36)<=signed(DIN_65_7)*signed(FMAP_37_65);
			MULT_66(36)<=signed(DIN_66_7)*signed(FMAP_37_66);
			MULT_67(36)<=signed(DIN_67_7)*signed(FMAP_37_67);
			MULT_68(36)<=signed(DIN_68_7)*signed(FMAP_37_68);
			MULT_69(36)<=signed(DIN_69_7)*signed(FMAP_37_69);
			MULT_70(36)<=signed(DIN_70_7)*signed(FMAP_37_70);
			MULT_71(36)<=signed(DIN_71_7)*signed(FMAP_37_71);
			MULT_72(36)<=signed(DIN_72_7)*signed(FMAP_37_72);
			MULT_73(36)<=signed(DIN_73_7)*signed(FMAP_37_73);
			MULT_74(36)<=signed(DIN_74_7)*signed(FMAP_37_74);
			MULT_75(36)<=signed(DIN_75_7)*signed(FMAP_37_75);
			MULT_76(36)<=signed(DIN_76_7)*signed(FMAP_37_76);
			MULT_77(36)<=signed(DIN_77_7)*signed(FMAP_37_77);
			MULT_78(36)<=signed(DIN_78_7)*signed(FMAP_37_78);
			MULT_79(36)<=signed(DIN_79_7)*signed(FMAP_37_79);
			MULT_80(36)<=signed(DIN_80_7)*signed(FMAP_37_80);
			MULT_81(36)<=signed(DIN_81_7)*signed(FMAP_37_81);
			MULT_82(36)<=signed(DIN_82_7)*signed(FMAP_37_82);
			MULT_83(36)<=signed(DIN_83_7)*signed(FMAP_37_83);
			MULT_84(36)<=signed(DIN_84_7)*signed(FMAP_37_84);
			MULT_85(36)<=signed(DIN_85_7)*signed(FMAP_37_85);
			MULT_86(36)<=signed(DIN_86_7)*signed(FMAP_37_86);
			MULT_87(36)<=signed(DIN_87_7)*signed(FMAP_37_87);
			MULT_88(36)<=signed(DIN_88_7)*signed(FMAP_37_88);
			MULT_89(36)<=signed(DIN_89_7)*signed(FMAP_37_89);
			MULT_90(36)<=signed(DIN_90_7)*signed(FMAP_37_90);
			MULT_91(36)<=signed(DIN_91_7)*signed(FMAP_37_91);
			MULT_92(36)<=signed(DIN_92_7)*signed(FMAP_37_92);
			MULT_93(36)<=signed(DIN_93_7)*signed(FMAP_37_93);
			MULT_94(36)<=signed(DIN_94_7)*signed(FMAP_37_94);
			MULT_95(36)<=signed(DIN_95_7)*signed(FMAP_37_95);
			MULT_96(36)<=signed(DIN_96_7)*signed(FMAP_37_96);
			MULT_97(36)<=signed(DIN_97_7)*signed(FMAP_37_97);
			MULT_98(36)<=signed(DIN_98_7)*signed(FMAP_37_98);
			MULT_99(36)<=signed(DIN_99_7)*signed(FMAP_37_99);
			MULT_100(36)<=signed(DIN_100_7)*signed(FMAP_37_100);
			MULT_101(36)<=signed(DIN_101_7)*signed(FMAP_37_101);
			MULT_102(36)<=signed(DIN_102_7)*signed(FMAP_37_102);
			MULT_103(36)<=signed(DIN_103_7)*signed(FMAP_37_103);
			MULT_104(36)<=signed(DIN_104_7)*signed(FMAP_37_104);
			MULT_105(36)<=signed(DIN_105_7)*signed(FMAP_37_105);
			MULT_106(36)<=signed(DIN_106_7)*signed(FMAP_37_106);
			MULT_107(36)<=signed(DIN_107_7)*signed(FMAP_37_107);
			MULT_108(36)<=signed(DIN_108_7)*signed(FMAP_37_108);
			MULT_109(36)<=signed(DIN_109_7)*signed(FMAP_37_109);
			MULT_110(36)<=signed(DIN_110_7)*signed(FMAP_37_110);
			MULT_111(36)<=signed(DIN_111_7)*signed(FMAP_37_111);
			MULT_112(36)<=signed(DIN_112_7)*signed(FMAP_37_112);
			MULT_113(36)<=signed(DIN_113_7)*signed(FMAP_37_113);
			MULT_114(36)<=signed(DIN_114_7)*signed(FMAP_37_114);
			MULT_115(36)<=signed(DIN_115_7)*signed(FMAP_37_115);
			MULT_116(36)<=signed(DIN_116_7)*signed(FMAP_37_116);
			MULT_117(36)<=signed(DIN_117_7)*signed(FMAP_37_117);
			MULT_118(36)<=signed(DIN_118_7)*signed(FMAP_37_118);
			MULT_119(36)<=signed(DIN_119_7)*signed(FMAP_37_119);
			MULT_120(36)<=signed(DIN_120_7)*signed(FMAP_37_120);

			MULT_1(37)<=signed(DIN_1_7)*signed(FMAP_38_1);
			MULT_2(37)<=signed(DIN_2_7)*signed(FMAP_38_2);
			MULT_3(37)<=signed(DIN_3_7)*signed(FMAP_38_3);
			MULT_4(37)<=signed(DIN_4_7)*signed(FMAP_38_4);
			MULT_5(37)<=signed(DIN_5_7)*signed(FMAP_38_5);
			MULT_6(37)<=signed(DIN_6_7)*signed(FMAP_38_6);
			MULT_7(37)<=signed(DIN_7_7)*signed(FMAP_38_7);
			MULT_8(37)<=signed(DIN_8_7)*signed(FMAP_38_8);
			MULT_9(37)<=signed(DIN_9_7)*signed(FMAP_38_9);
			MULT_10(37)<=signed(DIN_10_7)*signed(FMAP_38_10);
			MULT_11(37)<=signed(DIN_11_7)*signed(FMAP_38_11);
			MULT_12(37)<=signed(DIN_12_7)*signed(FMAP_38_12);
			MULT_13(37)<=signed(DIN_13_7)*signed(FMAP_38_13);
			MULT_14(37)<=signed(DIN_14_7)*signed(FMAP_38_14);
			MULT_15(37)<=signed(DIN_15_7)*signed(FMAP_38_15);
			MULT_16(37)<=signed(DIN_16_7)*signed(FMAP_38_16);
			MULT_17(37)<=signed(DIN_17_7)*signed(FMAP_38_17);
			MULT_18(37)<=signed(DIN_18_7)*signed(FMAP_38_18);
			MULT_19(37)<=signed(DIN_19_7)*signed(FMAP_38_19);
			MULT_20(37)<=signed(DIN_20_7)*signed(FMAP_38_20);
			MULT_21(37)<=signed(DIN_21_7)*signed(FMAP_38_21);
			MULT_22(37)<=signed(DIN_22_7)*signed(FMAP_38_22);
			MULT_23(37)<=signed(DIN_23_7)*signed(FMAP_38_23);
			MULT_24(37)<=signed(DIN_24_7)*signed(FMAP_38_24);
			MULT_25(37)<=signed(DIN_25_7)*signed(FMAP_38_25);
			MULT_26(37)<=signed(DIN_26_7)*signed(FMAP_38_26);
			MULT_27(37)<=signed(DIN_27_7)*signed(FMAP_38_27);
			MULT_28(37)<=signed(DIN_28_7)*signed(FMAP_38_28);
			MULT_29(37)<=signed(DIN_29_7)*signed(FMAP_38_29);
			MULT_30(37)<=signed(DIN_30_7)*signed(FMAP_38_30);
			MULT_31(37)<=signed(DIN_31_7)*signed(FMAP_38_31);
			MULT_32(37)<=signed(DIN_32_7)*signed(FMAP_38_32);
			MULT_33(37)<=signed(DIN_33_7)*signed(FMAP_38_33);
			MULT_34(37)<=signed(DIN_34_7)*signed(FMAP_38_34);
			MULT_35(37)<=signed(DIN_35_7)*signed(FMAP_38_35);
			MULT_36(37)<=signed(DIN_36_7)*signed(FMAP_38_36);
			MULT_37(37)<=signed(DIN_37_7)*signed(FMAP_38_37);
			MULT_38(37)<=signed(DIN_38_7)*signed(FMAP_38_38);
			MULT_39(37)<=signed(DIN_39_7)*signed(FMAP_38_39);
			MULT_40(37)<=signed(DIN_40_7)*signed(FMAP_38_40);
			MULT_41(37)<=signed(DIN_41_7)*signed(FMAP_38_41);
			MULT_42(37)<=signed(DIN_42_7)*signed(FMAP_38_42);
			MULT_43(37)<=signed(DIN_43_7)*signed(FMAP_38_43);
			MULT_44(37)<=signed(DIN_44_7)*signed(FMAP_38_44);
			MULT_45(37)<=signed(DIN_45_7)*signed(FMAP_38_45);
			MULT_46(37)<=signed(DIN_46_7)*signed(FMAP_38_46);
			MULT_47(37)<=signed(DIN_47_7)*signed(FMAP_38_47);
			MULT_48(37)<=signed(DIN_48_7)*signed(FMAP_38_48);
			MULT_49(37)<=signed(DIN_49_7)*signed(FMAP_38_49);
			MULT_50(37)<=signed(DIN_50_7)*signed(FMAP_38_50);
			MULT_51(37)<=signed(DIN_51_7)*signed(FMAP_38_51);
			MULT_52(37)<=signed(DIN_52_7)*signed(FMAP_38_52);
			MULT_53(37)<=signed(DIN_53_7)*signed(FMAP_38_53);
			MULT_54(37)<=signed(DIN_54_7)*signed(FMAP_38_54);
			MULT_55(37)<=signed(DIN_55_7)*signed(FMAP_38_55);
			MULT_56(37)<=signed(DIN_56_7)*signed(FMAP_38_56);
			MULT_57(37)<=signed(DIN_57_7)*signed(FMAP_38_57);
			MULT_58(37)<=signed(DIN_58_7)*signed(FMAP_38_58);
			MULT_59(37)<=signed(DIN_59_7)*signed(FMAP_38_59);
			MULT_60(37)<=signed(DIN_60_7)*signed(FMAP_38_60);
			MULT_61(37)<=signed(DIN_61_7)*signed(FMAP_38_61);
			MULT_62(37)<=signed(DIN_62_7)*signed(FMAP_38_62);
			MULT_63(37)<=signed(DIN_63_7)*signed(FMAP_38_63);
			MULT_64(37)<=signed(DIN_64_7)*signed(FMAP_38_64);
			MULT_65(37)<=signed(DIN_65_7)*signed(FMAP_38_65);
			MULT_66(37)<=signed(DIN_66_7)*signed(FMAP_38_66);
			MULT_67(37)<=signed(DIN_67_7)*signed(FMAP_38_67);
			MULT_68(37)<=signed(DIN_68_7)*signed(FMAP_38_68);
			MULT_69(37)<=signed(DIN_69_7)*signed(FMAP_38_69);
			MULT_70(37)<=signed(DIN_70_7)*signed(FMAP_38_70);
			MULT_71(37)<=signed(DIN_71_7)*signed(FMAP_38_71);
			MULT_72(37)<=signed(DIN_72_7)*signed(FMAP_38_72);
			MULT_73(37)<=signed(DIN_73_7)*signed(FMAP_38_73);
			MULT_74(37)<=signed(DIN_74_7)*signed(FMAP_38_74);
			MULT_75(37)<=signed(DIN_75_7)*signed(FMAP_38_75);
			MULT_76(37)<=signed(DIN_76_7)*signed(FMAP_38_76);
			MULT_77(37)<=signed(DIN_77_7)*signed(FMAP_38_77);
			MULT_78(37)<=signed(DIN_78_7)*signed(FMAP_38_78);
			MULT_79(37)<=signed(DIN_79_7)*signed(FMAP_38_79);
			MULT_80(37)<=signed(DIN_80_7)*signed(FMAP_38_80);
			MULT_81(37)<=signed(DIN_81_7)*signed(FMAP_38_81);
			MULT_82(37)<=signed(DIN_82_7)*signed(FMAP_38_82);
			MULT_83(37)<=signed(DIN_83_7)*signed(FMAP_38_83);
			MULT_84(37)<=signed(DIN_84_7)*signed(FMAP_38_84);
			MULT_85(37)<=signed(DIN_85_7)*signed(FMAP_38_85);
			MULT_86(37)<=signed(DIN_86_7)*signed(FMAP_38_86);
			MULT_87(37)<=signed(DIN_87_7)*signed(FMAP_38_87);
			MULT_88(37)<=signed(DIN_88_7)*signed(FMAP_38_88);
			MULT_89(37)<=signed(DIN_89_7)*signed(FMAP_38_89);
			MULT_90(37)<=signed(DIN_90_7)*signed(FMAP_38_90);
			MULT_91(37)<=signed(DIN_91_7)*signed(FMAP_38_91);
			MULT_92(37)<=signed(DIN_92_7)*signed(FMAP_38_92);
			MULT_93(37)<=signed(DIN_93_7)*signed(FMAP_38_93);
			MULT_94(37)<=signed(DIN_94_7)*signed(FMAP_38_94);
			MULT_95(37)<=signed(DIN_95_7)*signed(FMAP_38_95);
			MULT_96(37)<=signed(DIN_96_7)*signed(FMAP_38_96);
			MULT_97(37)<=signed(DIN_97_7)*signed(FMAP_38_97);
			MULT_98(37)<=signed(DIN_98_7)*signed(FMAP_38_98);
			MULT_99(37)<=signed(DIN_99_7)*signed(FMAP_38_99);
			MULT_100(37)<=signed(DIN_100_7)*signed(FMAP_38_100);
			MULT_101(37)<=signed(DIN_101_7)*signed(FMAP_38_101);
			MULT_102(37)<=signed(DIN_102_7)*signed(FMAP_38_102);
			MULT_103(37)<=signed(DIN_103_7)*signed(FMAP_38_103);
			MULT_104(37)<=signed(DIN_104_7)*signed(FMAP_38_104);
			MULT_105(37)<=signed(DIN_105_7)*signed(FMAP_38_105);
			MULT_106(37)<=signed(DIN_106_7)*signed(FMAP_38_106);
			MULT_107(37)<=signed(DIN_107_7)*signed(FMAP_38_107);
			MULT_108(37)<=signed(DIN_108_7)*signed(FMAP_38_108);
			MULT_109(37)<=signed(DIN_109_7)*signed(FMAP_38_109);
			MULT_110(37)<=signed(DIN_110_7)*signed(FMAP_38_110);
			MULT_111(37)<=signed(DIN_111_7)*signed(FMAP_38_111);
			MULT_112(37)<=signed(DIN_112_7)*signed(FMAP_38_112);
			MULT_113(37)<=signed(DIN_113_7)*signed(FMAP_38_113);
			MULT_114(37)<=signed(DIN_114_7)*signed(FMAP_38_114);
			MULT_115(37)<=signed(DIN_115_7)*signed(FMAP_38_115);
			MULT_116(37)<=signed(DIN_116_7)*signed(FMAP_38_116);
			MULT_117(37)<=signed(DIN_117_7)*signed(FMAP_38_117);
			MULT_118(37)<=signed(DIN_118_7)*signed(FMAP_38_118);
			MULT_119(37)<=signed(DIN_119_7)*signed(FMAP_38_119);
			MULT_120(37)<=signed(DIN_120_7)*signed(FMAP_38_120);

			MULT_1(38)<=signed(DIN_1_7)*signed(FMAP_39_1);
			MULT_2(38)<=signed(DIN_2_7)*signed(FMAP_39_2);
			MULT_3(38)<=signed(DIN_3_7)*signed(FMAP_39_3);
			MULT_4(38)<=signed(DIN_4_7)*signed(FMAP_39_4);
			MULT_5(38)<=signed(DIN_5_7)*signed(FMAP_39_5);
			MULT_6(38)<=signed(DIN_6_7)*signed(FMAP_39_6);
			MULT_7(38)<=signed(DIN_7_7)*signed(FMAP_39_7);
			MULT_8(38)<=signed(DIN_8_7)*signed(FMAP_39_8);
			MULT_9(38)<=signed(DIN_9_7)*signed(FMAP_39_9);
			MULT_10(38)<=signed(DIN_10_7)*signed(FMAP_39_10);
			MULT_11(38)<=signed(DIN_11_7)*signed(FMAP_39_11);
			MULT_12(38)<=signed(DIN_12_7)*signed(FMAP_39_12);
			MULT_13(38)<=signed(DIN_13_7)*signed(FMAP_39_13);
			MULT_14(38)<=signed(DIN_14_7)*signed(FMAP_39_14);
			MULT_15(38)<=signed(DIN_15_7)*signed(FMAP_39_15);
			MULT_16(38)<=signed(DIN_16_7)*signed(FMAP_39_16);
			MULT_17(38)<=signed(DIN_17_7)*signed(FMAP_39_17);
			MULT_18(38)<=signed(DIN_18_7)*signed(FMAP_39_18);
			MULT_19(38)<=signed(DIN_19_7)*signed(FMAP_39_19);
			MULT_20(38)<=signed(DIN_20_7)*signed(FMAP_39_20);
			MULT_21(38)<=signed(DIN_21_7)*signed(FMAP_39_21);
			MULT_22(38)<=signed(DIN_22_7)*signed(FMAP_39_22);
			MULT_23(38)<=signed(DIN_23_7)*signed(FMAP_39_23);
			MULT_24(38)<=signed(DIN_24_7)*signed(FMAP_39_24);
			MULT_25(38)<=signed(DIN_25_7)*signed(FMAP_39_25);
			MULT_26(38)<=signed(DIN_26_7)*signed(FMAP_39_26);
			MULT_27(38)<=signed(DIN_27_7)*signed(FMAP_39_27);
			MULT_28(38)<=signed(DIN_28_7)*signed(FMAP_39_28);
			MULT_29(38)<=signed(DIN_29_7)*signed(FMAP_39_29);
			MULT_30(38)<=signed(DIN_30_7)*signed(FMAP_39_30);
			MULT_31(38)<=signed(DIN_31_7)*signed(FMAP_39_31);
			MULT_32(38)<=signed(DIN_32_7)*signed(FMAP_39_32);
			MULT_33(38)<=signed(DIN_33_7)*signed(FMAP_39_33);
			MULT_34(38)<=signed(DIN_34_7)*signed(FMAP_39_34);
			MULT_35(38)<=signed(DIN_35_7)*signed(FMAP_39_35);
			MULT_36(38)<=signed(DIN_36_7)*signed(FMAP_39_36);
			MULT_37(38)<=signed(DIN_37_7)*signed(FMAP_39_37);
			MULT_38(38)<=signed(DIN_38_7)*signed(FMAP_39_38);
			MULT_39(38)<=signed(DIN_39_7)*signed(FMAP_39_39);
			MULT_40(38)<=signed(DIN_40_7)*signed(FMAP_39_40);
			MULT_41(38)<=signed(DIN_41_7)*signed(FMAP_39_41);
			MULT_42(38)<=signed(DIN_42_7)*signed(FMAP_39_42);
			MULT_43(38)<=signed(DIN_43_7)*signed(FMAP_39_43);
			MULT_44(38)<=signed(DIN_44_7)*signed(FMAP_39_44);
			MULT_45(38)<=signed(DIN_45_7)*signed(FMAP_39_45);
			MULT_46(38)<=signed(DIN_46_7)*signed(FMAP_39_46);
			MULT_47(38)<=signed(DIN_47_7)*signed(FMAP_39_47);
			MULT_48(38)<=signed(DIN_48_7)*signed(FMAP_39_48);
			MULT_49(38)<=signed(DIN_49_7)*signed(FMAP_39_49);
			MULT_50(38)<=signed(DIN_50_7)*signed(FMAP_39_50);
			MULT_51(38)<=signed(DIN_51_7)*signed(FMAP_39_51);
			MULT_52(38)<=signed(DIN_52_7)*signed(FMAP_39_52);
			MULT_53(38)<=signed(DIN_53_7)*signed(FMAP_39_53);
			MULT_54(38)<=signed(DIN_54_7)*signed(FMAP_39_54);
			MULT_55(38)<=signed(DIN_55_7)*signed(FMAP_39_55);
			MULT_56(38)<=signed(DIN_56_7)*signed(FMAP_39_56);
			MULT_57(38)<=signed(DIN_57_7)*signed(FMAP_39_57);
			MULT_58(38)<=signed(DIN_58_7)*signed(FMAP_39_58);
			MULT_59(38)<=signed(DIN_59_7)*signed(FMAP_39_59);
			MULT_60(38)<=signed(DIN_60_7)*signed(FMAP_39_60);
			MULT_61(38)<=signed(DIN_61_7)*signed(FMAP_39_61);
			MULT_62(38)<=signed(DIN_62_7)*signed(FMAP_39_62);
			MULT_63(38)<=signed(DIN_63_7)*signed(FMAP_39_63);
			MULT_64(38)<=signed(DIN_64_7)*signed(FMAP_39_64);
			MULT_65(38)<=signed(DIN_65_7)*signed(FMAP_39_65);
			MULT_66(38)<=signed(DIN_66_7)*signed(FMAP_39_66);
			MULT_67(38)<=signed(DIN_67_7)*signed(FMAP_39_67);
			MULT_68(38)<=signed(DIN_68_7)*signed(FMAP_39_68);
			MULT_69(38)<=signed(DIN_69_7)*signed(FMAP_39_69);
			MULT_70(38)<=signed(DIN_70_7)*signed(FMAP_39_70);
			MULT_71(38)<=signed(DIN_71_7)*signed(FMAP_39_71);
			MULT_72(38)<=signed(DIN_72_7)*signed(FMAP_39_72);
			MULT_73(38)<=signed(DIN_73_7)*signed(FMAP_39_73);
			MULT_74(38)<=signed(DIN_74_7)*signed(FMAP_39_74);
			MULT_75(38)<=signed(DIN_75_7)*signed(FMAP_39_75);
			MULT_76(38)<=signed(DIN_76_7)*signed(FMAP_39_76);
			MULT_77(38)<=signed(DIN_77_7)*signed(FMAP_39_77);
			MULT_78(38)<=signed(DIN_78_7)*signed(FMAP_39_78);
			MULT_79(38)<=signed(DIN_79_7)*signed(FMAP_39_79);
			MULT_80(38)<=signed(DIN_80_7)*signed(FMAP_39_80);
			MULT_81(38)<=signed(DIN_81_7)*signed(FMAP_39_81);
			MULT_82(38)<=signed(DIN_82_7)*signed(FMAP_39_82);
			MULT_83(38)<=signed(DIN_83_7)*signed(FMAP_39_83);
			MULT_84(38)<=signed(DIN_84_7)*signed(FMAP_39_84);
			MULT_85(38)<=signed(DIN_85_7)*signed(FMAP_39_85);
			MULT_86(38)<=signed(DIN_86_7)*signed(FMAP_39_86);
			MULT_87(38)<=signed(DIN_87_7)*signed(FMAP_39_87);
			MULT_88(38)<=signed(DIN_88_7)*signed(FMAP_39_88);
			MULT_89(38)<=signed(DIN_89_7)*signed(FMAP_39_89);
			MULT_90(38)<=signed(DIN_90_7)*signed(FMAP_39_90);
			MULT_91(38)<=signed(DIN_91_7)*signed(FMAP_39_91);
			MULT_92(38)<=signed(DIN_92_7)*signed(FMAP_39_92);
			MULT_93(38)<=signed(DIN_93_7)*signed(FMAP_39_93);
			MULT_94(38)<=signed(DIN_94_7)*signed(FMAP_39_94);
			MULT_95(38)<=signed(DIN_95_7)*signed(FMAP_39_95);
			MULT_96(38)<=signed(DIN_96_7)*signed(FMAP_39_96);
			MULT_97(38)<=signed(DIN_97_7)*signed(FMAP_39_97);
			MULT_98(38)<=signed(DIN_98_7)*signed(FMAP_39_98);
			MULT_99(38)<=signed(DIN_99_7)*signed(FMAP_39_99);
			MULT_100(38)<=signed(DIN_100_7)*signed(FMAP_39_100);
			MULT_101(38)<=signed(DIN_101_7)*signed(FMAP_39_101);
			MULT_102(38)<=signed(DIN_102_7)*signed(FMAP_39_102);
			MULT_103(38)<=signed(DIN_103_7)*signed(FMAP_39_103);
			MULT_104(38)<=signed(DIN_104_7)*signed(FMAP_39_104);
			MULT_105(38)<=signed(DIN_105_7)*signed(FMAP_39_105);
			MULT_106(38)<=signed(DIN_106_7)*signed(FMAP_39_106);
			MULT_107(38)<=signed(DIN_107_7)*signed(FMAP_39_107);
			MULT_108(38)<=signed(DIN_108_7)*signed(FMAP_39_108);
			MULT_109(38)<=signed(DIN_109_7)*signed(FMAP_39_109);
			MULT_110(38)<=signed(DIN_110_7)*signed(FMAP_39_110);
			MULT_111(38)<=signed(DIN_111_7)*signed(FMAP_39_111);
			MULT_112(38)<=signed(DIN_112_7)*signed(FMAP_39_112);
			MULT_113(38)<=signed(DIN_113_7)*signed(FMAP_39_113);
			MULT_114(38)<=signed(DIN_114_7)*signed(FMAP_39_114);
			MULT_115(38)<=signed(DIN_115_7)*signed(FMAP_39_115);
			MULT_116(38)<=signed(DIN_116_7)*signed(FMAP_39_116);
			MULT_117(38)<=signed(DIN_117_7)*signed(FMAP_39_117);
			MULT_118(38)<=signed(DIN_118_7)*signed(FMAP_39_118);
			MULT_119(38)<=signed(DIN_119_7)*signed(FMAP_39_119);
			MULT_120(38)<=signed(DIN_120_7)*signed(FMAP_39_120);

			MULT_1(39)<=signed(DIN_1_7)*signed(FMAP_40_1);
			MULT_2(39)<=signed(DIN_2_7)*signed(FMAP_40_2);
			MULT_3(39)<=signed(DIN_3_7)*signed(FMAP_40_3);
			MULT_4(39)<=signed(DIN_4_7)*signed(FMAP_40_4);
			MULT_5(39)<=signed(DIN_5_7)*signed(FMAP_40_5);
			MULT_6(39)<=signed(DIN_6_7)*signed(FMAP_40_6);
			MULT_7(39)<=signed(DIN_7_7)*signed(FMAP_40_7);
			MULT_8(39)<=signed(DIN_8_7)*signed(FMAP_40_8);
			MULT_9(39)<=signed(DIN_9_7)*signed(FMAP_40_9);
			MULT_10(39)<=signed(DIN_10_7)*signed(FMAP_40_10);
			MULT_11(39)<=signed(DIN_11_7)*signed(FMAP_40_11);
			MULT_12(39)<=signed(DIN_12_7)*signed(FMAP_40_12);
			MULT_13(39)<=signed(DIN_13_7)*signed(FMAP_40_13);
			MULT_14(39)<=signed(DIN_14_7)*signed(FMAP_40_14);
			MULT_15(39)<=signed(DIN_15_7)*signed(FMAP_40_15);
			MULT_16(39)<=signed(DIN_16_7)*signed(FMAP_40_16);
			MULT_17(39)<=signed(DIN_17_7)*signed(FMAP_40_17);
			MULT_18(39)<=signed(DIN_18_7)*signed(FMAP_40_18);
			MULT_19(39)<=signed(DIN_19_7)*signed(FMAP_40_19);
			MULT_20(39)<=signed(DIN_20_7)*signed(FMAP_40_20);
			MULT_21(39)<=signed(DIN_21_7)*signed(FMAP_40_21);
			MULT_22(39)<=signed(DIN_22_7)*signed(FMAP_40_22);
			MULT_23(39)<=signed(DIN_23_7)*signed(FMAP_40_23);
			MULT_24(39)<=signed(DIN_24_7)*signed(FMAP_40_24);
			MULT_25(39)<=signed(DIN_25_7)*signed(FMAP_40_25);
			MULT_26(39)<=signed(DIN_26_7)*signed(FMAP_40_26);
			MULT_27(39)<=signed(DIN_27_7)*signed(FMAP_40_27);
			MULT_28(39)<=signed(DIN_28_7)*signed(FMAP_40_28);
			MULT_29(39)<=signed(DIN_29_7)*signed(FMAP_40_29);
			MULT_30(39)<=signed(DIN_30_7)*signed(FMAP_40_30);
			MULT_31(39)<=signed(DIN_31_7)*signed(FMAP_40_31);
			MULT_32(39)<=signed(DIN_32_7)*signed(FMAP_40_32);
			MULT_33(39)<=signed(DIN_33_7)*signed(FMAP_40_33);
			MULT_34(39)<=signed(DIN_34_7)*signed(FMAP_40_34);
			MULT_35(39)<=signed(DIN_35_7)*signed(FMAP_40_35);
			MULT_36(39)<=signed(DIN_36_7)*signed(FMAP_40_36);
			MULT_37(39)<=signed(DIN_37_7)*signed(FMAP_40_37);
			MULT_38(39)<=signed(DIN_38_7)*signed(FMAP_40_38);
			MULT_39(39)<=signed(DIN_39_7)*signed(FMAP_40_39);
			MULT_40(39)<=signed(DIN_40_7)*signed(FMAP_40_40);
			MULT_41(39)<=signed(DIN_41_7)*signed(FMAP_40_41);
			MULT_42(39)<=signed(DIN_42_7)*signed(FMAP_40_42);
			MULT_43(39)<=signed(DIN_43_7)*signed(FMAP_40_43);
			MULT_44(39)<=signed(DIN_44_7)*signed(FMAP_40_44);
			MULT_45(39)<=signed(DIN_45_7)*signed(FMAP_40_45);
			MULT_46(39)<=signed(DIN_46_7)*signed(FMAP_40_46);
			MULT_47(39)<=signed(DIN_47_7)*signed(FMAP_40_47);
			MULT_48(39)<=signed(DIN_48_7)*signed(FMAP_40_48);
			MULT_49(39)<=signed(DIN_49_7)*signed(FMAP_40_49);
			MULT_50(39)<=signed(DIN_50_7)*signed(FMAP_40_50);
			MULT_51(39)<=signed(DIN_51_7)*signed(FMAP_40_51);
			MULT_52(39)<=signed(DIN_52_7)*signed(FMAP_40_52);
			MULT_53(39)<=signed(DIN_53_7)*signed(FMAP_40_53);
			MULT_54(39)<=signed(DIN_54_7)*signed(FMAP_40_54);
			MULT_55(39)<=signed(DIN_55_7)*signed(FMAP_40_55);
			MULT_56(39)<=signed(DIN_56_7)*signed(FMAP_40_56);
			MULT_57(39)<=signed(DIN_57_7)*signed(FMAP_40_57);
			MULT_58(39)<=signed(DIN_58_7)*signed(FMAP_40_58);
			MULT_59(39)<=signed(DIN_59_7)*signed(FMAP_40_59);
			MULT_60(39)<=signed(DIN_60_7)*signed(FMAP_40_60);
			MULT_61(39)<=signed(DIN_61_7)*signed(FMAP_40_61);
			MULT_62(39)<=signed(DIN_62_7)*signed(FMAP_40_62);
			MULT_63(39)<=signed(DIN_63_7)*signed(FMAP_40_63);
			MULT_64(39)<=signed(DIN_64_7)*signed(FMAP_40_64);
			MULT_65(39)<=signed(DIN_65_7)*signed(FMAP_40_65);
			MULT_66(39)<=signed(DIN_66_7)*signed(FMAP_40_66);
			MULT_67(39)<=signed(DIN_67_7)*signed(FMAP_40_67);
			MULT_68(39)<=signed(DIN_68_7)*signed(FMAP_40_68);
			MULT_69(39)<=signed(DIN_69_7)*signed(FMAP_40_69);
			MULT_70(39)<=signed(DIN_70_7)*signed(FMAP_40_70);
			MULT_71(39)<=signed(DIN_71_7)*signed(FMAP_40_71);
			MULT_72(39)<=signed(DIN_72_7)*signed(FMAP_40_72);
			MULT_73(39)<=signed(DIN_73_7)*signed(FMAP_40_73);
			MULT_74(39)<=signed(DIN_74_7)*signed(FMAP_40_74);
			MULT_75(39)<=signed(DIN_75_7)*signed(FMAP_40_75);
			MULT_76(39)<=signed(DIN_76_7)*signed(FMAP_40_76);
			MULT_77(39)<=signed(DIN_77_7)*signed(FMAP_40_77);
			MULT_78(39)<=signed(DIN_78_7)*signed(FMAP_40_78);
			MULT_79(39)<=signed(DIN_79_7)*signed(FMAP_40_79);
			MULT_80(39)<=signed(DIN_80_7)*signed(FMAP_40_80);
			MULT_81(39)<=signed(DIN_81_7)*signed(FMAP_40_81);
			MULT_82(39)<=signed(DIN_82_7)*signed(FMAP_40_82);
			MULT_83(39)<=signed(DIN_83_7)*signed(FMAP_40_83);
			MULT_84(39)<=signed(DIN_84_7)*signed(FMAP_40_84);
			MULT_85(39)<=signed(DIN_85_7)*signed(FMAP_40_85);
			MULT_86(39)<=signed(DIN_86_7)*signed(FMAP_40_86);
			MULT_87(39)<=signed(DIN_87_7)*signed(FMAP_40_87);
			MULT_88(39)<=signed(DIN_88_7)*signed(FMAP_40_88);
			MULT_89(39)<=signed(DIN_89_7)*signed(FMAP_40_89);
			MULT_90(39)<=signed(DIN_90_7)*signed(FMAP_40_90);
			MULT_91(39)<=signed(DIN_91_7)*signed(FMAP_40_91);
			MULT_92(39)<=signed(DIN_92_7)*signed(FMAP_40_92);
			MULT_93(39)<=signed(DIN_93_7)*signed(FMAP_40_93);
			MULT_94(39)<=signed(DIN_94_7)*signed(FMAP_40_94);
			MULT_95(39)<=signed(DIN_95_7)*signed(FMAP_40_95);
			MULT_96(39)<=signed(DIN_96_7)*signed(FMAP_40_96);
			MULT_97(39)<=signed(DIN_97_7)*signed(FMAP_40_97);
			MULT_98(39)<=signed(DIN_98_7)*signed(FMAP_40_98);
			MULT_99(39)<=signed(DIN_99_7)*signed(FMAP_40_99);
			MULT_100(39)<=signed(DIN_100_7)*signed(FMAP_40_100);
			MULT_101(39)<=signed(DIN_101_7)*signed(FMAP_40_101);
			MULT_102(39)<=signed(DIN_102_7)*signed(FMAP_40_102);
			MULT_103(39)<=signed(DIN_103_7)*signed(FMAP_40_103);
			MULT_104(39)<=signed(DIN_104_7)*signed(FMAP_40_104);
			MULT_105(39)<=signed(DIN_105_7)*signed(FMAP_40_105);
			MULT_106(39)<=signed(DIN_106_7)*signed(FMAP_40_106);
			MULT_107(39)<=signed(DIN_107_7)*signed(FMAP_40_107);
			MULT_108(39)<=signed(DIN_108_7)*signed(FMAP_40_108);
			MULT_109(39)<=signed(DIN_109_7)*signed(FMAP_40_109);
			MULT_110(39)<=signed(DIN_110_7)*signed(FMAP_40_110);
			MULT_111(39)<=signed(DIN_111_7)*signed(FMAP_40_111);
			MULT_112(39)<=signed(DIN_112_7)*signed(FMAP_40_112);
			MULT_113(39)<=signed(DIN_113_7)*signed(FMAP_40_113);
			MULT_114(39)<=signed(DIN_114_7)*signed(FMAP_40_114);
			MULT_115(39)<=signed(DIN_115_7)*signed(FMAP_40_115);
			MULT_116(39)<=signed(DIN_116_7)*signed(FMAP_40_116);
			MULT_117(39)<=signed(DIN_117_7)*signed(FMAP_40_117);
			MULT_118(39)<=signed(DIN_118_7)*signed(FMAP_40_118);
			MULT_119(39)<=signed(DIN_119_7)*signed(FMAP_40_119);
			MULT_120(39)<=signed(DIN_120_7)*signed(FMAP_40_120);

			MULT_1(40)<=signed(DIN_1_7)*signed(FMAP_41_1);
			MULT_2(40)<=signed(DIN_2_7)*signed(FMAP_41_2);
			MULT_3(40)<=signed(DIN_3_7)*signed(FMAP_41_3);
			MULT_4(40)<=signed(DIN_4_7)*signed(FMAP_41_4);
			MULT_5(40)<=signed(DIN_5_7)*signed(FMAP_41_5);
			MULT_6(40)<=signed(DIN_6_7)*signed(FMAP_41_6);
			MULT_7(40)<=signed(DIN_7_7)*signed(FMAP_41_7);
			MULT_8(40)<=signed(DIN_8_7)*signed(FMAP_41_8);
			MULT_9(40)<=signed(DIN_9_7)*signed(FMAP_41_9);
			MULT_10(40)<=signed(DIN_10_7)*signed(FMAP_41_10);
			MULT_11(40)<=signed(DIN_11_7)*signed(FMAP_41_11);
			MULT_12(40)<=signed(DIN_12_7)*signed(FMAP_41_12);
			MULT_13(40)<=signed(DIN_13_7)*signed(FMAP_41_13);
			MULT_14(40)<=signed(DIN_14_7)*signed(FMAP_41_14);
			MULT_15(40)<=signed(DIN_15_7)*signed(FMAP_41_15);
			MULT_16(40)<=signed(DIN_16_7)*signed(FMAP_41_16);
			MULT_17(40)<=signed(DIN_17_7)*signed(FMAP_41_17);
			MULT_18(40)<=signed(DIN_18_7)*signed(FMAP_41_18);
			MULT_19(40)<=signed(DIN_19_7)*signed(FMAP_41_19);
			MULT_20(40)<=signed(DIN_20_7)*signed(FMAP_41_20);
			MULT_21(40)<=signed(DIN_21_7)*signed(FMAP_41_21);
			MULT_22(40)<=signed(DIN_22_7)*signed(FMAP_41_22);
			MULT_23(40)<=signed(DIN_23_7)*signed(FMAP_41_23);
			MULT_24(40)<=signed(DIN_24_7)*signed(FMAP_41_24);
			MULT_25(40)<=signed(DIN_25_7)*signed(FMAP_41_25);
			MULT_26(40)<=signed(DIN_26_7)*signed(FMAP_41_26);
			MULT_27(40)<=signed(DIN_27_7)*signed(FMAP_41_27);
			MULT_28(40)<=signed(DIN_28_7)*signed(FMAP_41_28);
			MULT_29(40)<=signed(DIN_29_7)*signed(FMAP_41_29);
			MULT_30(40)<=signed(DIN_30_7)*signed(FMAP_41_30);
			MULT_31(40)<=signed(DIN_31_7)*signed(FMAP_41_31);
			MULT_32(40)<=signed(DIN_32_7)*signed(FMAP_41_32);
			MULT_33(40)<=signed(DIN_33_7)*signed(FMAP_41_33);
			MULT_34(40)<=signed(DIN_34_7)*signed(FMAP_41_34);
			MULT_35(40)<=signed(DIN_35_7)*signed(FMAP_41_35);
			MULT_36(40)<=signed(DIN_36_7)*signed(FMAP_41_36);
			MULT_37(40)<=signed(DIN_37_7)*signed(FMAP_41_37);
			MULT_38(40)<=signed(DIN_38_7)*signed(FMAP_41_38);
			MULT_39(40)<=signed(DIN_39_7)*signed(FMAP_41_39);
			MULT_40(40)<=signed(DIN_40_7)*signed(FMAP_41_40);
			MULT_41(40)<=signed(DIN_41_7)*signed(FMAP_41_41);
			MULT_42(40)<=signed(DIN_42_7)*signed(FMAP_41_42);
			MULT_43(40)<=signed(DIN_43_7)*signed(FMAP_41_43);
			MULT_44(40)<=signed(DIN_44_7)*signed(FMAP_41_44);
			MULT_45(40)<=signed(DIN_45_7)*signed(FMAP_41_45);
			MULT_46(40)<=signed(DIN_46_7)*signed(FMAP_41_46);
			MULT_47(40)<=signed(DIN_47_7)*signed(FMAP_41_47);
			MULT_48(40)<=signed(DIN_48_7)*signed(FMAP_41_48);
			MULT_49(40)<=signed(DIN_49_7)*signed(FMAP_41_49);
			MULT_50(40)<=signed(DIN_50_7)*signed(FMAP_41_50);
			MULT_51(40)<=signed(DIN_51_7)*signed(FMAP_41_51);
			MULT_52(40)<=signed(DIN_52_7)*signed(FMAP_41_52);
			MULT_53(40)<=signed(DIN_53_7)*signed(FMAP_41_53);
			MULT_54(40)<=signed(DIN_54_7)*signed(FMAP_41_54);
			MULT_55(40)<=signed(DIN_55_7)*signed(FMAP_41_55);
			MULT_56(40)<=signed(DIN_56_7)*signed(FMAP_41_56);
			MULT_57(40)<=signed(DIN_57_7)*signed(FMAP_41_57);
			MULT_58(40)<=signed(DIN_58_7)*signed(FMAP_41_58);
			MULT_59(40)<=signed(DIN_59_7)*signed(FMAP_41_59);
			MULT_60(40)<=signed(DIN_60_7)*signed(FMAP_41_60);
			MULT_61(40)<=signed(DIN_61_7)*signed(FMAP_41_61);
			MULT_62(40)<=signed(DIN_62_7)*signed(FMAP_41_62);
			MULT_63(40)<=signed(DIN_63_7)*signed(FMAP_41_63);
			MULT_64(40)<=signed(DIN_64_7)*signed(FMAP_41_64);
			MULT_65(40)<=signed(DIN_65_7)*signed(FMAP_41_65);
			MULT_66(40)<=signed(DIN_66_7)*signed(FMAP_41_66);
			MULT_67(40)<=signed(DIN_67_7)*signed(FMAP_41_67);
			MULT_68(40)<=signed(DIN_68_7)*signed(FMAP_41_68);
			MULT_69(40)<=signed(DIN_69_7)*signed(FMAP_41_69);
			MULT_70(40)<=signed(DIN_70_7)*signed(FMAP_41_70);
			MULT_71(40)<=signed(DIN_71_7)*signed(FMAP_41_71);
			MULT_72(40)<=signed(DIN_72_7)*signed(FMAP_41_72);
			MULT_73(40)<=signed(DIN_73_7)*signed(FMAP_41_73);
			MULT_74(40)<=signed(DIN_74_7)*signed(FMAP_41_74);
			MULT_75(40)<=signed(DIN_75_7)*signed(FMAP_41_75);
			MULT_76(40)<=signed(DIN_76_7)*signed(FMAP_41_76);
			MULT_77(40)<=signed(DIN_77_7)*signed(FMAP_41_77);
			MULT_78(40)<=signed(DIN_78_7)*signed(FMAP_41_78);
			MULT_79(40)<=signed(DIN_79_7)*signed(FMAP_41_79);
			MULT_80(40)<=signed(DIN_80_7)*signed(FMAP_41_80);
			MULT_81(40)<=signed(DIN_81_7)*signed(FMAP_41_81);
			MULT_82(40)<=signed(DIN_82_7)*signed(FMAP_41_82);
			MULT_83(40)<=signed(DIN_83_7)*signed(FMAP_41_83);
			MULT_84(40)<=signed(DIN_84_7)*signed(FMAP_41_84);
			MULT_85(40)<=signed(DIN_85_7)*signed(FMAP_41_85);
			MULT_86(40)<=signed(DIN_86_7)*signed(FMAP_41_86);
			MULT_87(40)<=signed(DIN_87_7)*signed(FMAP_41_87);
			MULT_88(40)<=signed(DIN_88_7)*signed(FMAP_41_88);
			MULT_89(40)<=signed(DIN_89_7)*signed(FMAP_41_89);
			MULT_90(40)<=signed(DIN_90_7)*signed(FMAP_41_90);
			MULT_91(40)<=signed(DIN_91_7)*signed(FMAP_41_91);
			MULT_92(40)<=signed(DIN_92_7)*signed(FMAP_41_92);
			MULT_93(40)<=signed(DIN_93_7)*signed(FMAP_41_93);
			MULT_94(40)<=signed(DIN_94_7)*signed(FMAP_41_94);
			MULT_95(40)<=signed(DIN_95_7)*signed(FMAP_41_95);
			MULT_96(40)<=signed(DIN_96_7)*signed(FMAP_41_96);
			MULT_97(40)<=signed(DIN_97_7)*signed(FMAP_41_97);
			MULT_98(40)<=signed(DIN_98_7)*signed(FMAP_41_98);
			MULT_99(40)<=signed(DIN_99_7)*signed(FMAP_41_99);
			MULT_100(40)<=signed(DIN_100_7)*signed(FMAP_41_100);
			MULT_101(40)<=signed(DIN_101_7)*signed(FMAP_41_101);
			MULT_102(40)<=signed(DIN_102_7)*signed(FMAP_41_102);
			MULT_103(40)<=signed(DIN_103_7)*signed(FMAP_41_103);
			MULT_104(40)<=signed(DIN_104_7)*signed(FMAP_41_104);
			MULT_105(40)<=signed(DIN_105_7)*signed(FMAP_41_105);
			MULT_106(40)<=signed(DIN_106_7)*signed(FMAP_41_106);
			MULT_107(40)<=signed(DIN_107_7)*signed(FMAP_41_107);
			MULT_108(40)<=signed(DIN_108_7)*signed(FMAP_41_108);
			MULT_109(40)<=signed(DIN_109_7)*signed(FMAP_41_109);
			MULT_110(40)<=signed(DIN_110_7)*signed(FMAP_41_110);
			MULT_111(40)<=signed(DIN_111_7)*signed(FMAP_41_111);
			MULT_112(40)<=signed(DIN_112_7)*signed(FMAP_41_112);
			MULT_113(40)<=signed(DIN_113_7)*signed(FMAP_41_113);
			MULT_114(40)<=signed(DIN_114_7)*signed(FMAP_41_114);
			MULT_115(40)<=signed(DIN_115_7)*signed(FMAP_41_115);
			MULT_116(40)<=signed(DIN_116_7)*signed(FMAP_41_116);
			MULT_117(40)<=signed(DIN_117_7)*signed(FMAP_41_117);
			MULT_118(40)<=signed(DIN_118_7)*signed(FMAP_41_118);
			MULT_119(40)<=signed(DIN_119_7)*signed(FMAP_41_119);
			MULT_120(40)<=signed(DIN_120_7)*signed(FMAP_41_120);

			MULT_1(41)<=signed(DIN_1_7)*signed(FMAP_42_1);
			MULT_2(41)<=signed(DIN_2_7)*signed(FMAP_42_2);
			MULT_3(41)<=signed(DIN_3_7)*signed(FMAP_42_3);
			MULT_4(41)<=signed(DIN_4_7)*signed(FMAP_42_4);
			MULT_5(41)<=signed(DIN_5_7)*signed(FMAP_42_5);
			MULT_6(41)<=signed(DIN_6_7)*signed(FMAP_42_6);
			MULT_7(41)<=signed(DIN_7_7)*signed(FMAP_42_7);
			MULT_8(41)<=signed(DIN_8_7)*signed(FMAP_42_8);
			MULT_9(41)<=signed(DIN_9_7)*signed(FMAP_42_9);
			MULT_10(41)<=signed(DIN_10_7)*signed(FMAP_42_10);
			MULT_11(41)<=signed(DIN_11_7)*signed(FMAP_42_11);
			MULT_12(41)<=signed(DIN_12_7)*signed(FMAP_42_12);
			MULT_13(41)<=signed(DIN_13_7)*signed(FMAP_42_13);
			MULT_14(41)<=signed(DIN_14_7)*signed(FMAP_42_14);
			MULT_15(41)<=signed(DIN_15_7)*signed(FMAP_42_15);
			MULT_16(41)<=signed(DIN_16_7)*signed(FMAP_42_16);
			MULT_17(41)<=signed(DIN_17_7)*signed(FMAP_42_17);
			MULT_18(41)<=signed(DIN_18_7)*signed(FMAP_42_18);
			MULT_19(41)<=signed(DIN_19_7)*signed(FMAP_42_19);
			MULT_20(41)<=signed(DIN_20_7)*signed(FMAP_42_20);
			MULT_21(41)<=signed(DIN_21_7)*signed(FMAP_42_21);
			MULT_22(41)<=signed(DIN_22_7)*signed(FMAP_42_22);
			MULT_23(41)<=signed(DIN_23_7)*signed(FMAP_42_23);
			MULT_24(41)<=signed(DIN_24_7)*signed(FMAP_42_24);
			MULT_25(41)<=signed(DIN_25_7)*signed(FMAP_42_25);
			MULT_26(41)<=signed(DIN_26_7)*signed(FMAP_42_26);
			MULT_27(41)<=signed(DIN_27_7)*signed(FMAP_42_27);
			MULT_28(41)<=signed(DIN_28_7)*signed(FMAP_42_28);
			MULT_29(41)<=signed(DIN_29_7)*signed(FMAP_42_29);
			MULT_30(41)<=signed(DIN_30_7)*signed(FMAP_42_30);
			MULT_31(41)<=signed(DIN_31_7)*signed(FMAP_42_31);
			MULT_32(41)<=signed(DIN_32_7)*signed(FMAP_42_32);
			MULT_33(41)<=signed(DIN_33_7)*signed(FMAP_42_33);
			MULT_34(41)<=signed(DIN_34_7)*signed(FMAP_42_34);
			MULT_35(41)<=signed(DIN_35_7)*signed(FMAP_42_35);
			MULT_36(41)<=signed(DIN_36_7)*signed(FMAP_42_36);
			MULT_37(41)<=signed(DIN_37_7)*signed(FMAP_42_37);
			MULT_38(41)<=signed(DIN_38_7)*signed(FMAP_42_38);
			MULT_39(41)<=signed(DIN_39_7)*signed(FMAP_42_39);
			MULT_40(41)<=signed(DIN_40_7)*signed(FMAP_42_40);
			MULT_41(41)<=signed(DIN_41_7)*signed(FMAP_42_41);
			MULT_42(41)<=signed(DIN_42_7)*signed(FMAP_42_42);
			MULT_43(41)<=signed(DIN_43_7)*signed(FMAP_42_43);
			MULT_44(41)<=signed(DIN_44_7)*signed(FMAP_42_44);
			MULT_45(41)<=signed(DIN_45_7)*signed(FMAP_42_45);
			MULT_46(41)<=signed(DIN_46_7)*signed(FMAP_42_46);
			MULT_47(41)<=signed(DIN_47_7)*signed(FMAP_42_47);
			MULT_48(41)<=signed(DIN_48_7)*signed(FMAP_42_48);
			MULT_49(41)<=signed(DIN_49_7)*signed(FMAP_42_49);
			MULT_50(41)<=signed(DIN_50_7)*signed(FMAP_42_50);
			MULT_51(41)<=signed(DIN_51_7)*signed(FMAP_42_51);
			MULT_52(41)<=signed(DIN_52_7)*signed(FMAP_42_52);
			MULT_53(41)<=signed(DIN_53_7)*signed(FMAP_42_53);
			MULT_54(41)<=signed(DIN_54_7)*signed(FMAP_42_54);
			MULT_55(41)<=signed(DIN_55_7)*signed(FMAP_42_55);
			MULT_56(41)<=signed(DIN_56_7)*signed(FMAP_42_56);
			MULT_57(41)<=signed(DIN_57_7)*signed(FMAP_42_57);
			MULT_58(41)<=signed(DIN_58_7)*signed(FMAP_42_58);
			MULT_59(41)<=signed(DIN_59_7)*signed(FMAP_42_59);
			MULT_60(41)<=signed(DIN_60_7)*signed(FMAP_42_60);
			MULT_61(41)<=signed(DIN_61_7)*signed(FMAP_42_61);
			MULT_62(41)<=signed(DIN_62_7)*signed(FMAP_42_62);
			MULT_63(41)<=signed(DIN_63_7)*signed(FMAP_42_63);
			MULT_64(41)<=signed(DIN_64_7)*signed(FMAP_42_64);
			MULT_65(41)<=signed(DIN_65_7)*signed(FMAP_42_65);
			MULT_66(41)<=signed(DIN_66_7)*signed(FMAP_42_66);
			MULT_67(41)<=signed(DIN_67_7)*signed(FMAP_42_67);
			MULT_68(41)<=signed(DIN_68_7)*signed(FMAP_42_68);
			MULT_69(41)<=signed(DIN_69_7)*signed(FMAP_42_69);
			MULT_70(41)<=signed(DIN_70_7)*signed(FMAP_42_70);
			MULT_71(41)<=signed(DIN_71_7)*signed(FMAP_42_71);
			MULT_72(41)<=signed(DIN_72_7)*signed(FMAP_42_72);
			MULT_73(41)<=signed(DIN_73_7)*signed(FMAP_42_73);
			MULT_74(41)<=signed(DIN_74_7)*signed(FMAP_42_74);
			MULT_75(41)<=signed(DIN_75_7)*signed(FMAP_42_75);
			MULT_76(41)<=signed(DIN_76_7)*signed(FMAP_42_76);
			MULT_77(41)<=signed(DIN_77_7)*signed(FMAP_42_77);
			MULT_78(41)<=signed(DIN_78_7)*signed(FMAP_42_78);
			MULT_79(41)<=signed(DIN_79_7)*signed(FMAP_42_79);
			MULT_80(41)<=signed(DIN_80_7)*signed(FMAP_42_80);
			MULT_81(41)<=signed(DIN_81_7)*signed(FMAP_42_81);
			MULT_82(41)<=signed(DIN_82_7)*signed(FMAP_42_82);
			MULT_83(41)<=signed(DIN_83_7)*signed(FMAP_42_83);
			MULT_84(41)<=signed(DIN_84_7)*signed(FMAP_42_84);
			MULT_85(41)<=signed(DIN_85_7)*signed(FMAP_42_85);
			MULT_86(41)<=signed(DIN_86_7)*signed(FMAP_42_86);
			MULT_87(41)<=signed(DIN_87_7)*signed(FMAP_42_87);
			MULT_88(41)<=signed(DIN_88_7)*signed(FMAP_42_88);
			MULT_89(41)<=signed(DIN_89_7)*signed(FMAP_42_89);
			MULT_90(41)<=signed(DIN_90_7)*signed(FMAP_42_90);
			MULT_91(41)<=signed(DIN_91_7)*signed(FMAP_42_91);
			MULT_92(41)<=signed(DIN_92_7)*signed(FMAP_42_92);
			MULT_93(41)<=signed(DIN_93_7)*signed(FMAP_42_93);
			MULT_94(41)<=signed(DIN_94_7)*signed(FMAP_42_94);
			MULT_95(41)<=signed(DIN_95_7)*signed(FMAP_42_95);
			MULT_96(41)<=signed(DIN_96_7)*signed(FMAP_42_96);
			MULT_97(41)<=signed(DIN_97_7)*signed(FMAP_42_97);
			MULT_98(41)<=signed(DIN_98_7)*signed(FMAP_42_98);
			MULT_99(41)<=signed(DIN_99_7)*signed(FMAP_42_99);
			MULT_100(41)<=signed(DIN_100_7)*signed(FMAP_42_100);
			MULT_101(41)<=signed(DIN_101_7)*signed(FMAP_42_101);
			MULT_102(41)<=signed(DIN_102_7)*signed(FMAP_42_102);
			MULT_103(41)<=signed(DIN_103_7)*signed(FMAP_42_103);
			MULT_104(41)<=signed(DIN_104_7)*signed(FMAP_42_104);
			MULT_105(41)<=signed(DIN_105_7)*signed(FMAP_42_105);
			MULT_106(41)<=signed(DIN_106_7)*signed(FMAP_42_106);
			MULT_107(41)<=signed(DIN_107_7)*signed(FMAP_42_107);
			MULT_108(41)<=signed(DIN_108_7)*signed(FMAP_42_108);
			MULT_109(41)<=signed(DIN_109_7)*signed(FMAP_42_109);
			MULT_110(41)<=signed(DIN_110_7)*signed(FMAP_42_110);
			MULT_111(41)<=signed(DIN_111_7)*signed(FMAP_42_111);
			MULT_112(41)<=signed(DIN_112_7)*signed(FMAP_42_112);
			MULT_113(41)<=signed(DIN_113_7)*signed(FMAP_42_113);
			MULT_114(41)<=signed(DIN_114_7)*signed(FMAP_42_114);
			MULT_115(41)<=signed(DIN_115_7)*signed(FMAP_42_115);
			MULT_116(41)<=signed(DIN_116_7)*signed(FMAP_42_116);
			MULT_117(41)<=signed(DIN_117_7)*signed(FMAP_42_117);
			MULT_118(41)<=signed(DIN_118_7)*signed(FMAP_42_118);
			MULT_119(41)<=signed(DIN_119_7)*signed(FMAP_42_119);
			MULT_120(41)<=signed(DIN_120_7)*signed(FMAP_42_120);

			MULT_1(42)<=signed(DIN_1_7)*signed(FMAP_43_1);
			MULT_2(42)<=signed(DIN_2_7)*signed(FMAP_43_2);
			MULT_3(42)<=signed(DIN_3_7)*signed(FMAP_43_3);
			MULT_4(42)<=signed(DIN_4_7)*signed(FMAP_43_4);
			MULT_5(42)<=signed(DIN_5_7)*signed(FMAP_43_5);
			MULT_6(42)<=signed(DIN_6_7)*signed(FMAP_43_6);
			MULT_7(42)<=signed(DIN_7_7)*signed(FMAP_43_7);
			MULT_8(42)<=signed(DIN_8_7)*signed(FMAP_43_8);
			MULT_9(42)<=signed(DIN_9_7)*signed(FMAP_43_9);
			MULT_10(42)<=signed(DIN_10_7)*signed(FMAP_43_10);
			MULT_11(42)<=signed(DIN_11_7)*signed(FMAP_43_11);
			MULT_12(42)<=signed(DIN_12_7)*signed(FMAP_43_12);
			MULT_13(42)<=signed(DIN_13_7)*signed(FMAP_43_13);
			MULT_14(42)<=signed(DIN_14_7)*signed(FMAP_43_14);
			MULT_15(42)<=signed(DIN_15_7)*signed(FMAP_43_15);
			MULT_16(42)<=signed(DIN_16_7)*signed(FMAP_43_16);
			MULT_17(42)<=signed(DIN_17_7)*signed(FMAP_43_17);
			MULT_18(42)<=signed(DIN_18_7)*signed(FMAP_43_18);
			MULT_19(42)<=signed(DIN_19_7)*signed(FMAP_43_19);
			MULT_20(42)<=signed(DIN_20_7)*signed(FMAP_43_20);
			MULT_21(42)<=signed(DIN_21_7)*signed(FMAP_43_21);
			MULT_22(42)<=signed(DIN_22_7)*signed(FMAP_43_22);
			MULT_23(42)<=signed(DIN_23_7)*signed(FMAP_43_23);
			MULT_24(42)<=signed(DIN_24_7)*signed(FMAP_43_24);
			MULT_25(42)<=signed(DIN_25_7)*signed(FMAP_43_25);
			MULT_26(42)<=signed(DIN_26_7)*signed(FMAP_43_26);
			MULT_27(42)<=signed(DIN_27_7)*signed(FMAP_43_27);
			MULT_28(42)<=signed(DIN_28_7)*signed(FMAP_43_28);
			MULT_29(42)<=signed(DIN_29_7)*signed(FMAP_43_29);
			MULT_30(42)<=signed(DIN_30_7)*signed(FMAP_43_30);
			MULT_31(42)<=signed(DIN_31_7)*signed(FMAP_43_31);
			MULT_32(42)<=signed(DIN_32_7)*signed(FMAP_43_32);
			MULT_33(42)<=signed(DIN_33_7)*signed(FMAP_43_33);
			MULT_34(42)<=signed(DIN_34_7)*signed(FMAP_43_34);
			MULT_35(42)<=signed(DIN_35_7)*signed(FMAP_43_35);
			MULT_36(42)<=signed(DIN_36_7)*signed(FMAP_43_36);
			MULT_37(42)<=signed(DIN_37_7)*signed(FMAP_43_37);
			MULT_38(42)<=signed(DIN_38_7)*signed(FMAP_43_38);
			MULT_39(42)<=signed(DIN_39_7)*signed(FMAP_43_39);
			MULT_40(42)<=signed(DIN_40_7)*signed(FMAP_43_40);
			MULT_41(42)<=signed(DIN_41_7)*signed(FMAP_43_41);
			MULT_42(42)<=signed(DIN_42_7)*signed(FMAP_43_42);
			MULT_43(42)<=signed(DIN_43_7)*signed(FMAP_43_43);
			MULT_44(42)<=signed(DIN_44_7)*signed(FMAP_43_44);
			MULT_45(42)<=signed(DIN_45_7)*signed(FMAP_43_45);
			MULT_46(42)<=signed(DIN_46_7)*signed(FMAP_43_46);
			MULT_47(42)<=signed(DIN_47_7)*signed(FMAP_43_47);
			MULT_48(42)<=signed(DIN_48_7)*signed(FMAP_43_48);
			MULT_49(42)<=signed(DIN_49_7)*signed(FMAP_43_49);
			MULT_50(42)<=signed(DIN_50_7)*signed(FMAP_43_50);
			MULT_51(42)<=signed(DIN_51_7)*signed(FMAP_43_51);
			MULT_52(42)<=signed(DIN_52_7)*signed(FMAP_43_52);
			MULT_53(42)<=signed(DIN_53_7)*signed(FMAP_43_53);
			MULT_54(42)<=signed(DIN_54_7)*signed(FMAP_43_54);
			MULT_55(42)<=signed(DIN_55_7)*signed(FMAP_43_55);
			MULT_56(42)<=signed(DIN_56_7)*signed(FMAP_43_56);
			MULT_57(42)<=signed(DIN_57_7)*signed(FMAP_43_57);
			MULT_58(42)<=signed(DIN_58_7)*signed(FMAP_43_58);
			MULT_59(42)<=signed(DIN_59_7)*signed(FMAP_43_59);
			MULT_60(42)<=signed(DIN_60_7)*signed(FMAP_43_60);
			MULT_61(42)<=signed(DIN_61_7)*signed(FMAP_43_61);
			MULT_62(42)<=signed(DIN_62_7)*signed(FMAP_43_62);
			MULT_63(42)<=signed(DIN_63_7)*signed(FMAP_43_63);
			MULT_64(42)<=signed(DIN_64_7)*signed(FMAP_43_64);
			MULT_65(42)<=signed(DIN_65_7)*signed(FMAP_43_65);
			MULT_66(42)<=signed(DIN_66_7)*signed(FMAP_43_66);
			MULT_67(42)<=signed(DIN_67_7)*signed(FMAP_43_67);
			MULT_68(42)<=signed(DIN_68_7)*signed(FMAP_43_68);
			MULT_69(42)<=signed(DIN_69_7)*signed(FMAP_43_69);
			MULT_70(42)<=signed(DIN_70_7)*signed(FMAP_43_70);
			MULT_71(42)<=signed(DIN_71_7)*signed(FMAP_43_71);
			MULT_72(42)<=signed(DIN_72_7)*signed(FMAP_43_72);
			MULT_73(42)<=signed(DIN_73_7)*signed(FMAP_43_73);
			MULT_74(42)<=signed(DIN_74_7)*signed(FMAP_43_74);
			MULT_75(42)<=signed(DIN_75_7)*signed(FMAP_43_75);
			MULT_76(42)<=signed(DIN_76_7)*signed(FMAP_43_76);
			MULT_77(42)<=signed(DIN_77_7)*signed(FMAP_43_77);
			MULT_78(42)<=signed(DIN_78_7)*signed(FMAP_43_78);
			MULT_79(42)<=signed(DIN_79_7)*signed(FMAP_43_79);
			MULT_80(42)<=signed(DIN_80_7)*signed(FMAP_43_80);
			MULT_81(42)<=signed(DIN_81_7)*signed(FMAP_43_81);
			MULT_82(42)<=signed(DIN_82_7)*signed(FMAP_43_82);
			MULT_83(42)<=signed(DIN_83_7)*signed(FMAP_43_83);
			MULT_84(42)<=signed(DIN_84_7)*signed(FMAP_43_84);
			MULT_85(42)<=signed(DIN_85_7)*signed(FMAP_43_85);
			MULT_86(42)<=signed(DIN_86_7)*signed(FMAP_43_86);
			MULT_87(42)<=signed(DIN_87_7)*signed(FMAP_43_87);
			MULT_88(42)<=signed(DIN_88_7)*signed(FMAP_43_88);
			MULT_89(42)<=signed(DIN_89_7)*signed(FMAP_43_89);
			MULT_90(42)<=signed(DIN_90_7)*signed(FMAP_43_90);
			MULT_91(42)<=signed(DIN_91_7)*signed(FMAP_43_91);
			MULT_92(42)<=signed(DIN_92_7)*signed(FMAP_43_92);
			MULT_93(42)<=signed(DIN_93_7)*signed(FMAP_43_93);
			MULT_94(42)<=signed(DIN_94_7)*signed(FMAP_43_94);
			MULT_95(42)<=signed(DIN_95_7)*signed(FMAP_43_95);
			MULT_96(42)<=signed(DIN_96_7)*signed(FMAP_43_96);
			MULT_97(42)<=signed(DIN_97_7)*signed(FMAP_43_97);
			MULT_98(42)<=signed(DIN_98_7)*signed(FMAP_43_98);
			MULT_99(42)<=signed(DIN_99_7)*signed(FMAP_43_99);
			MULT_100(42)<=signed(DIN_100_7)*signed(FMAP_43_100);
			MULT_101(42)<=signed(DIN_101_7)*signed(FMAP_43_101);
			MULT_102(42)<=signed(DIN_102_7)*signed(FMAP_43_102);
			MULT_103(42)<=signed(DIN_103_7)*signed(FMAP_43_103);
			MULT_104(42)<=signed(DIN_104_7)*signed(FMAP_43_104);
			MULT_105(42)<=signed(DIN_105_7)*signed(FMAP_43_105);
			MULT_106(42)<=signed(DIN_106_7)*signed(FMAP_43_106);
			MULT_107(42)<=signed(DIN_107_7)*signed(FMAP_43_107);
			MULT_108(42)<=signed(DIN_108_7)*signed(FMAP_43_108);
			MULT_109(42)<=signed(DIN_109_7)*signed(FMAP_43_109);
			MULT_110(42)<=signed(DIN_110_7)*signed(FMAP_43_110);
			MULT_111(42)<=signed(DIN_111_7)*signed(FMAP_43_111);
			MULT_112(42)<=signed(DIN_112_7)*signed(FMAP_43_112);
			MULT_113(42)<=signed(DIN_113_7)*signed(FMAP_43_113);
			MULT_114(42)<=signed(DIN_114_7)*signed(FMAP_43_114);
			MULT_115(42)<=signed(DIN_115_7)*signed(FMAP_43_115);
			MULT_116(42)<=signed(DIN_116_7)*signed(FMAP_43_116);
			MULT_117(42)<=signed(DIN_117_7)*signed(FMAP_43_117);
			MULT_118(42)<=signed(DIN_118_7)*signed(FMAP_43_118);
			MULT_119(42)<=signed(DIN_119_7)*signed(FMAP_43_119);
			MULT_120(42)<=signed(DIN_120_7)*signed(FMAP_43_120);

			MULT_1(43)<=signed(DIN_1_7)*signed(FMAP_44_1);
			MULT_2(43)<=signed(DIN_2_7)*signed(FMAP_44_2);
			MULT_3(43)<=signed(DIN_3_7)*signed(FMAP_44_3);
			MULT_4(43)<=signed(DIN_4_7)*signed(FMAP_44_4);
			MULT_5(43)<=signed(DIN_5_7)*signed(FMAP_44_5);
			MULT_6(43)<=signed(DIN_6_7)*signed(FMAP_44_6);
			MULT_7(43)<=signed(DIN_7_7)*signed(FMAP_44_7);
			MULT_8(43)<=signed(DIN_8_7)*signed(FMAP_44_8);
			MULT_9(43)<=signed(DIN_9_7)*signed(FMAP_44_9);
			MULT_10(43)<=signed(DIN_10_7)*signed(FMAP_44_10);
			MULT_11(43)<=signed(DIN_11_7)*signed(FMAP_44_11);
			MULT_12(43)<=signed(DIN_12_7)*signed(FMAP_44_12);
			MULT_13(43)<=signed(DIN_13_7)*signed(FMAP_44_13);
			MULT_14(43)<=signed(DIN_14_7)*signed(FMAP_44_14);
			MULT_15(43)<=signed(DIN_15_7)*signed(FMAP_44_15);
			MULT_16(43)<=signed(DIN_16_7)*signed(FMAP_44_16);
			MULT_17(43)<=signed(DIN_17_7)*signed(FMAP_44_17);
			MULT_18(43)<=signed(DIN_18_7)*signed(FMAP_44_18);
			MULT_19(43)<=signed(DIN_19_7)*signed(FMAP_44_19);
			MULT_20(43)<=signed(DIN_20_7)*signed(FMAP_44_20);
			MULT_21(43)<=signed(DIN_21_7)*signed(FMAP_44_21);
			MULT_22(43)<=signed(DIN_22_7)*signed(FMAP_44_22);
			MULT_23(43)<=signed(DIN_23_7)*signed(FMAP_44_23);
			MULT_24(43)<=signed(DIN_24_7)*signed(FMAP_44_24);
			MULT_25(43)<=signed(DIN_25_7)*signed(FMAP_44_25);
			MULT_26(43)<=signed(DIN_26_7)*signed(FMAP_44_26);
			MULT_27(43)<=signed(DIN_27_7)*signed(FMAP_44_27);
			MULT_28(43)<=signed(DIN_28_7)*signed(FMAP_44_28);
			MULT_29(43)<=signed(DIN_29_7)*signed(FMAP_44_29);
			MULT_30(43)<=signed(DIN_30_7)*signed(FMAP_44_30);
			MULT_31(43)<=signed(DIN_31_7)*signed(FMAP_44_31);
			MULT_32(43)<=signed(DIN_32_7)*signed(FMAP_44_32);
			MULT_33(43)<=signed(DIN_33_7)*signed(FMAP_44_33);
			MULT_34(43)<=signed(DIN_34_7)*signed(FMAP_44_34);
			MULT_35(43)<=signed(DIN_35_7)*signed(FMAP_44_35);
			MULT_36(43)<=signed(DIN_36_7)*signed(FMAP_44_36);
			MULT_37(43)<=signed(DIN_37_7)*signed(FMAP_44_37);
			MULT_38(43)<=signed(DIN_38_7)*signed(FMAP_44_38);
			MULT_39(43)<=signed(DIN_39_7)*signed(FMAP_44_39);
			MULT_40(43)<=signed(DIN_40_7)*signed(FMAP_44_40);
			MULT_41(43)<=signed(DIN_41_7)*signed(FMAP_44_41);
			MULT_42(43)<=signed(DIN_42_7)*signed(FMAP_44_42);
			MULT_43(43)<=signed(DIN_43_7)*signed(FMAP_44_43);
			MULT_44(43)<=signed(DIN_44_7)*signed(FMAP_44_44);
			MULT_45(43)<=signed(DIN_45_7)*signed(FMAP_44_45);
			MULT_46(43)<=signed(DIN_46_7)*signed(FMAP_44_46);
			MULT_47(43)<=signed(DIN_47_7)*signed(FMAP_44_47);
			MULT_48(43)<=signed(DIN_48_7)*signed(FMAP_44_48);
			MULT_49(43)<=signed(DIN_49_7)*signed(FMAP_44_49);
			MULT_50(43)<=signed(DIN_50_7)*signed(FMAP_44_50);
			MULT_51(43)<=signed(DIN_51_7)*signed(FMAP_44_51);
			MULT_52(43)<=signed(DIN_52_7)*signed(FMAP_44_52);
			MULT_53(43)<=signed(DIN_53_7)*signed(FMAP_44_53);
			MULT_54(43)<=signed(DIN_54_7)*signed(FMAP_44_54);
			MULT_55(43)<=signed(DIN_55_7)*signed(FMAP_44_55);
			MULT_56(43)<=signed(DIN_56_7)*signed(FMAP_44_56);
			MULT_57(43)<=signed(DIN_57_7)*signed(FMAP_44_57);
			MULT_58(43)<=signed(DIN_58_7)*signed(FMAP_44_58);
			MULT_59(43)<=signed(DIN_59_7)*signed(FMAP_44_59);
			MULT_60(43)<=signed(DIN_60_7)*signed(FMAP_44_60);
			MULT_61(43)<=signed(DIN_61_7)*signed(FMAP_44_61);
			MULT_62(43)<=signed(DIN_62_7)*signed(FMAP_44_62);
			MULT_63(43)<=signed(DIN_63_7)*signed(FMAP_44_63);
			MULT_64(43)<=signed(DIN_64_7)*signed(FMAP_44_64);
			MULT_65(43)<=signed(DIN_65_7)*signed(FMAP_44_65);
			MULT_66(43)<=signed(DIN_66_7)*signed(FMAP_44_66);
			MULT_67(43)<=signed(DIN_67_7)*signed(FMAP_44_67);
			MULT_68(43)<=signed(DIN_68_7)*signed(FMAP_44_68);
			MULT_69(43)<=signed(DIN_69_7)*signed(FMAP_44_69);
			MULT_70(43)<=signed(DIN_70_7)*signed(FMAP_44_70);
			MULT_71(43)<=signed(DIN_71_7)*signed(FMAP_44_71);
			MULT_72(43)<=signed(DIN_72_7)*signed(FMAP_44_72);
			MULT_73(43)<=signed(DIN_73_7)*signed(FMAP_44_73);
			MULT_74(43)<=signed(DIN_74_7)*signed(FMAP_44_74);
			MULT_75(43)<=signed(DIN_75_7)*signed(FMAP_44_75);
			MULT_76(43)<=signed(DIN_76_7)*signed(FMAP_44_76);
			MULT_77(43)<=signed(DIN_77_7)*signed(FMAP_44_77);
			MULT_78(43)<=signed(DIN_78_7)*signed(FMAP_44_78);
			MULT_79(43)<=signed(DIN_79_7)*signed(FMAP_44_79);
			MULT_80(43)<=signed(DIN_80_7)*signed(FMAP_44_80);
			MULT_81(43)<=signed(DIN_81_7)*signed(FMAP_44_81);
			MULT_82(43)<=signed(DIN_82_7)*signed(FMAP_44_82);
			MULT_83(43)<=signed(DIN_83_7)*signed(FMAP_44_83);
			MULT_84(43)<=signed(DIN_84_7)*signed(FMAP_44_84);
			MULT_85(43)<=signed(DIN_85_7)*signed(FMAP_44_85);
			MULT_86(43)<=signed(DIN_86_7)*signed(FMAP_44_86);
			MULT_87(43)<=signed(DIN_87_7)*signed(FMAP_44_87);
			MULT_88(43)<=signed(DIN_88_7)*signed(FMAP_44_88);
			MULT_89(43)<=signed(DIN_89_7)*signed(FMAP_44_89);
			MULT_90(43)<=signed(DIN_90_7)*signed(FMAP_44_90);
			MULT_91(43)<=signed(DIN_91_7)*signed(FMAP_44_91);
			MULT_92(43)<=signed(DIN_92_7)*signed(FMAP_44_92);
			MULT_93(43)<=signed(DIN_93_7)*signed(FMAP_44_93);
			MULT_94(43)<=signed(DIN_94_7)*signed(FMAP_44_94);
			MULT_95(43)<=signed(DIN_95_7)*signed(FMAP_44_95);
			MULT_96(43)<=signed(DIN_96_7)*signed(FMAP_44_96);
			MULT_97(43)<=signed(DIN_97_7)*signed(FMAP_44_97);
			MULT_98(43)<=signed(DIN_98_7)*signed(FMAP_44_98);
			MULT_99(43)<=signed(DIN_99_7)*signed(FMAP_44_99);
			MULT_100(43)<=signed(DIN_100_7)*signed(FMAP_44_100);
			MULT_101(43)<=signed(DIN_101_7)*signed(FMAP_44_101);
			MULT_102(43)<=signed(DIN_102_7)*signed(FMAP_44_102);
			MULT_103(43)<=signed(DIN_103_7)*signed(FMAP_44_103);
			MULT_104(43)<=signed(DIN_104_7)*signed(FMAP_44_104);
			MULT_105(43)<=signed(DIN_105_7)*signed(FMAP_44_105);
			MULT_106(43)<=signed(DIN_106_7)*signed(FMAP_44_106);
			MULT_107(43)<=signed(DIN_107_7)*signed(FMAP_44_107);
			MULT_108(43)<=signed(DIN_108_7)*signed(FMAP_44_108);
			MULT_109(43)<=signed(DIN_109_7)*signed(FMAP_44_109);
			MULT_110(43)<=signed(DIN_110_7)*signed(FMAP_44_110);
			MULT_111(43)<=signed(DIN_111_7)*signed(FMAP_44_111);
			MULT_112(43)<=signed(DIN_112_7)*signed(FMAP_44_112);
			MULT_113(43)<=signed(DIN_113_7)*signed(FMAP_44_113);
			MULT_114(43)<=signed(DIN_114_7)*signed(FMAP_44_114);
			MULT_115(43)<=signed(DIN_115_7)*signed(FMAP_44_115);
			MULT_116(43)<=signed(DIN_116_7)*signed(FMAP_44_116);
			MULT_117(43)<=signed(DIN_117_7)*signed(FMAP_44_117);
			MULT_118(43)<=signed(DIN_118_7)*signed(FMAP_44_118);
			MULT_119(43)<=signed(DIN_119_7)*signed(FMAP_44_119);
			MULT_120(43)<=signed(DIN_120_7)*signed(FMAP_44_120);

			MULT_1(44)<=signed(DIN_1_7)*signed(FMAP_45_1);
			MULT_2(44)<=signed(DIN_2_7)*signed(FMAP_45_2);
			MULT_3(44)<=signed(DIN_3_7)*signed(FMAP_45_3);
			MULT_4(44)<=signed(DIN_4_7)*signed(FMAP_45_4);
			MULT_5(44)<=signed(DIN_5_7)*signed(FMAP_45_5);
			MULT_6(44)<=signed(DIN_6_7)*signed(FMAP_45_6);
			MULT_7(44)<=signed(DIN_7_7)*signed(FMAP_45_7);
			MULT_8(44)<=signed(DIN_8_7)*signed(FMAP_45_8);
			MULT_9(44)<=signed(DIN_9_7)*signed(FMAP_45_9);
			MULT_10(44)<=signed(DIN_10_7)*signed(FMAP_45_10);
			MULT_11(44)<=signed(DIN_11_7)*signed(FMAP_45_11);
			MULT_12(44)<=signed(DIN_12_7)*signed(FMAP_45_12);
			MULT_13(44)<=signed(DIN_13_7)*signed(FMAP_45_13);
			MULT_14(44)<=signed(DIN_14_7)*signed(FMAP_45_14);
			MULT_15(44)<=signed(DIN_15_7)*signed(FMAP_45_15);
			MULT_16(44)<=signed(DIN_16_7)*signed(FMAP_45_16);
			MULT_17(44)<=signed(DIN_17_7)*signed(FMAP_45_17);
			MULT_18(44)<=signed(DIN_18_7)*signed(FMAP_45_18);
			MULT_19(44)<=signed(DIN_19_7)*signed(FMAP_45_19);
			MULT_20(44)<=signed(DIN_20_7)*signed(FMAP_45_20);
			MULT_21(44)<=signed(DIN_21_7)*signed(FMAP_45_21);
			MULT_22(44)<=signed(DIN_22_7)*signed(FMAP_45_22);
			MULT_23(44)<=signed(DIN_23_7)*signed(FMAP_45_23);
			MULT_24(44)<=signed(DIN_24_7)*signed(FMAP_45_24);
			MULT_25(44)<=signed(DIN_25_7)*signed(FMAP_45_25);
			MULT_26(44)<=signed(DIN_26_7)*signed(FMAP_45_26);
			MULT_27(44)<=signed(DIN_27_7)*signed(FMAP_45_27);
			MULT_28(44)<=signed(DIN_28_7)*signed(FMAP_45_28);
			MULT_29(44)<=signed(DIN_29_7)*signed(FMAP_45_29);
			MULT_30(44)<=signed(DIN_30_7)*signed(FMAP_45_30);
			MULT_31(44)<=signed(DIN_31_7)*signed(FMAP_45_31);
			MULT_32(44)<=signed(DIN_32_7)*signed(FMAP_45_32);
			MULT_33(44)<=signed(DIN_33_7)*signed(FMAP_45_33);
			MULT_34(44)<=signed(DIN_34_7)*signed(FMAP_45_34);
			MULT_35(44)<=signed(DIN_35_7)*signed(FMAP_45_35);
			MULT_36(44)<=signed(DIN_36_7)*signed(FMAP_45_36);
			MULT_37(44)<=signed(DIN_37_7)*signed(FMAP_45_37);
			MULT_38(44)<=signed(DIN_38_7)*signed(FMAP_45_38);
			MULT_39(44)<=signed(DIN_39_7)*signed(FMAP_45_39);
			MULT_40(44)<=signed(DIN_40_7)*signed(FMAP_45_40);
			MULT_41(44)<=signed(DIN_41_7)*signed(FMAP_45_41);
			MULT_42(44)<=signed(DIN_42_7)*signed(FMAP_45_42);
			MULT_43(44)<=signed(DIN_43_7)*signed(FMAP_45_43);
			MULT_44(44)<=signed(DIN_44_7)*signed(FMAP_45_44);
			MULT_45(44)<=signed(DIN_45_7)*signed(FMAP_45_45);
			MULT_46(44)<=signed(DIN_46_7)*signed(FMAP_45_46);
			MULT_47(44)<=signed(DIN_47_7)*signed(FMAP_45_47);
			MULT_48(44)<=signed(DIN_48_7)*signed(FMAP_45_48);
			MULT_49(44)<=signed(DIN_49_7)*signed(FMAP_45_49);
			MULT_50(44)<=signed(DIN_50_7)*signed(FMAP_45_50);
			MULT_51(44)<=signed(DIN_51_7)*signed(FMAP_45_51);
			MULT_52(44)<=signed(DIN_52_7)*signed(FMAP_45_52);
			MULT_53(44)<=signed(DIN_53_7)*signed(FMAP_45_53);
			MULT_54(44)<=signed(DIN_54_7)*signed(FMAP_45_54);
			MULT_55(44)<=signed(DIN_55_7)*signed(FMAP_45_55);
			MULT_56(44)<=signed(DIN_56_7)*signed(FMAP_45_56);
			MULT_57(44)<=signed(DIN_57_7)*signed(FMAP_45_57);
			MULT_58(44)<=signed(DIN_58_7)*signed(FMAP_45_58);
			MULT_59(44)<=signed(DIN_59_7)*signed(FMAP_45_59);
			MULT_60(44)<=signed(DIN_60_7)*signed(FMAP_45_60);
			MULT_61(44)<=signed(DIN_61_7)*signed(FMAP_45_61);
			MULT_62(44)<=signed(DIN_62_7)*signed(FMAP_45_62);
			MULT_63(44)<=signed(DIN_63_7)*signed(FMAP_45_63);
			MULT_64(44)<=signed(DIN_64_7)*signed(FMAP_45_64);
			MULT_65(44)<=signed(DIN_65_7)*signed(FMAP_45_65);
			MULT_66(44)<=signed(DIN_66_7)*signed(FMAP_45_66);
			MULT_67(44)<=signed(DIN_67_7)*signed(FMAP_45_67);
			MULT_68(44)<=signed(DIN_68_7)*signed(FMAP_45_68);
			MULT_69(44)<=signed(DIN_69_7)*signed(FMAP_45_69);
			MULT_70(44)<=signed(DIN_70_7)*signed(FMAP_45_70);
			MULT_71(44)<=signed(DIN_71_7)*signed(FMAP_45_71);
			MULT_72(44)<=signed(DIN_72_7)*signed(FMAP_45_72);
			MULT_73(44)<=signed(DIN_73_7)*signed(FMAP_45_73);
			MULT_74(44)<=signed(DIN_74_7)*signed(FMAP_45_74);
			MULT_75(44)<=signed(DIN_75_7)*signed(FMAP_45_75);
			MULT_76(44)<=signed(DIN_76_7)*signed(FMAP_45_76);
			MULT_77(44)<=signed(DIN_77_7)*signed(FMAP_45_77);
			MULT_78(44)<=signed(DIN_78_7)*signed(FMAP_45_78);
			MULT_79(44)<=signed(DIN_79_7)*signed(FMAP_45_79);
			MULT_80(44)<=signed(DIN_80_7)*signed(FMAP_45_80);
			MULT_81(44)<=signed(DIN_81_7)*signed(FMAP_45_81);
			MULT_82(44)<=signed(DIN_82_7)*signed(FMAP_45_82);
			MULT_83(44)<=signed(DIN_83_7)*signed(FMAP_45_83);
			MULT_84(44)<=signed(DIN_84_7)*signed(FMAP_45_84);
			MULT_85(44)<=signed(DIN_85_7)*signed(FMAP_45_85);
			MULT_86(44)<=signed(DIN_86_7)*signed(FMAP_45_86);
			MULT_87(44)<=signed(DIN_87_7)*signed(FMAP_45_87);
			MULT_88(44)<=signed(DIN_88_7)*signed(FMAP_45_88);
			MULT_89(44)<=signed(DIN_89_7)*signed(FMAP_45_89);
			MULT_90(44)<=signed(DIN_90_7)*signed(FMAP_45_90);
			MULT_91(44)<=signed(DIN_91_7)*signed(FMAP_45_91);
			MULT_92(44)<=signed(DIN_92_7)*signed(FMAP_45_92);
			MULT_93(44)<=signed(DIN_93_7)*signed(FMAP_45_93);
			MULT_94(44)<=signed(DIN_94_7)*signed(FMAP_45_94);
			MULT_95(44)<=signed(DIN_95_7)*signed(FMAP_45_95);
			MULT_96(44)<=signed(DIN_96_7)*signed(FMAP_45_96);
			MULT_97(44)<=signed(DIN_97_7)*signed(FMAP_45_97);
			MULT_98(44)<=signed(DIN_98_7)*signed(FMAP_45_98);
			MULT_99(44)<=signed(DIN_99_7)*signed(FMAP_45_99);
			MULT_100(44)<=signed(DIN_100_7)*signed(FMAP_45_100);
			MULT_101(44)<=signed(DIN_101_7)*signed(FMAP_45_101);
			MULT_102(44)<=signed(DIN_102_7)*signed(FMAP_45_102);
			MULT_103(44)<=signed(DIN_103_7)*signed(FMAP_45_103);
			MULT_104(44)<=signed(DIN_104_7)*signed(FMAP_45_104);
			MULT_105(44)<=signed(DIN_105_7)*signed(FMAP_45_105);
			MULT_106(44)<=signed(DIN_106_7)*signed(FMAP_45_106);
			MULT_107(44)<=signed(DIN_107_7)*signed(FMAP_45_107);
			MULT_108(44)<=signed(DIN_108_7)*signed(FMAP_45_108);
			MULT_109(44)<=signed(DIN_109_7)*signed(FMAP_45_109);
			MULT_110(44)<=signed(DIN_110_7)*signed(FMAP_45_110);
			MULT_111(44)<=signed(DIN_111_7)*signed(FMAP_45_111);
			MULT_112(44)<=signed(DIN_112_7)*signed(FMAP_45_112);
			MULT_113(44)<=signed(DIN_113_7)*signed(FMAP_45_113);
			MULT_114(44)<=signed(DIN_114_7)*signed(FMAP_45_114);
			MULT_115(44)<=signed(DIN_115_7)*signed(FMAP_45_115);
			MULT_116(44)<=signed(DIN_116_7)*signed(FMAP_45_116);
			MULT_117(44)<=signed(DIN_117_7)*signed(FMAP_45_117);
			MULT_118(44)<=signed(DIN_118_7)*signed(FMAP_45_118);
			MULT_119(44)<=signed(DIN_119_7)*signed(FMAP_45_119);
			MULT_120(44)<=signed(DIN_120_7)*signed(FMAP_45_120);

			MULT_1(45)<=signed(DIN_1_7)*signed(FMAP_46_1);
			MULT_2(45)<=signed(DIN_2_7)*signed(FMAP_46_2);
			MULT_3(45)<=signed(DIN_3_7)*signed(FMAP_46_3);
			MULT_4(45)<=signed(DIN_4_7)*signed(FMAP_46_4);
			MULT_5(45)<=signed(DIN_5_7)*signed(FMAP_46_5);
			MULT_6(45)<=signed(DIN_6_7)*signed(FMAP_46_6);
			MULT_7(45)<=signed(DIN_7_7)*signed(FMAP_46_7);
			MULT_8(45)<=signed(DIN_8_7)*signed(FMAP_46_8);
			MULT_9(45)<=signed(DIN_9_7)*signed(FMAP_46_9);
			MULT_10(45)<=signed(DIN_10_7)*signed(FMAP_46_10);
			MULT_11(45)<=signed(DIN_11_7)*signed(FMAP_46_11);
			MULT_12(45)<=signed(DIN_12_7)*signed(FMAP_46_12);
			MULT_13(45)<=signed(DIN_13_7)*signed(FMAP_46_13);
			MULT_14(45)<=signed(DIN_14_7)*signed(FMAP_46_14);
			MULT_15(45)<=signed(DIN_15_7)*signed(FMAP_46_15);
			MULT_16(45)<=signed(DIN_16_7)*signed(FMAP_46_16);
			MULT_17(45)<=signed(DIN_17_7)*signed(FMAP_46_17);
			MULT_18(45)<=signed(DIN_18_7)*signed(FMAP_46_18);
			MULT_19(45)<=signed(DIN_19_7)*signed(FMAP_46_19);
			MULT_20(45)<=signed(DIN_20_7)*signed(FMAP_46_20);
			MULT_21(45)<=signed(DIN_21_7)*signed(FMAP_46_21);
			MULT_22(45)<=signed(DIN_22_7)*signed(FMAP_46_22);
			MULT_23(45)<=signed(DIN_23_7)*signed(FMAP_46_23);
			MULT_24(45)<=signed(DIN_24_7)*signed(FMAP_46_24);
			MULT_25(45)<=signed(DIN_25_7)*signed(FMAP_46_25);
			MULT_26(45)<=signed(DIN_26_7)*signed(FMAP_46_26);
			MULT_27(45)<=signed(DIN_27_7)*signed(FMAP_46_27);
			MULT_28(45)<=signed(DIN_28_7)*signed(FMAP_46_28);
			MULT_29(45)<=signed(DIN_29_7)*signed(FMAP_46_29);
			MULT_30(45)<=signed(DIN_30_7)*signed(FMAP_46_30);
			MULT_31(45)<=signed(DIN_31_7)*signed(FMAP_46_31);
			MULT_32(45)<=signed(DIN_32_7)*signed(FMAP_46_32);
			MULT_33(45)<=signed(DIN_33_7)*signed(FMAP_46_33);
			MULT_34(45)<=signed(DIN_34_7)*signed(FMAP_46_34);
			MULT_35(45)<=signed(DIN_35_7)*signed(FMAP_46_35);
			MULT_36(45)<=signed(DIN_36_7)*signed(FMAP_46_36);
			MULT_37(45)<=signed(DIN_37_7)*signed(FMAP_46_37);
			MULT_38(45)<=signed(DIN_38_7)*signed(FMAP_46_38);
			MULT_39(45)<=signed(DIN_39_7)*signed(FMAP_46_39);
			MULT_40(45)<=signed(DIN_40_7)*signed(FMAP_46_40);
			MULT_41(45)<=signed(DIN_41_7)*signed(FMAP_46_41);
			MULT_42(45)<=signed(DIN_42_7)*signed(FMAP_46_42);
			MULT_43(45)<=signed(DIN_43_7)*signed(FMAP_46_43);
			MULT_44(45)<=signed(DIN_44_7)*signed(FMAP_46_44);
			MULT_45(45)<=signed(DIN_45_7)*signed(FMAP_46_45);
			MULT_46(45)<=signed(DIN_46_7)*signed(FMAP_46_46);
			MULT_47(45)<=signed(DIN_47_7)*signed(FMAP_46_47);
			MULT_48(45)<=signed(DIN_48_7)*signed(FMAP_46_48);
			MULT_49(45)<=signed(DIN_49_7)*signed(FMAP_46_49);
			MULT_50(45)<=signed(DIN_50_7)*signed(FMAP_46_50);
			MULT_51(45)<=signed(DIN_51_7)*signed(FMAP_46_51);
			MULT_52(45)<=signed(DIN_52_7)*signed(FMAP_46_52);
			MULT_53(45)<=signed(DIN_53_7)*signed(FMAP_46_53);
			MULT_54(45)<=signed(DIN_54_7)*signed(FMAP_46_54);
			MULT_55(45)<=signed(DIN_55_7)*signed(FMAP_46_55);
			MULT_56(45)<=signed(DIN_56_7)*signed(FMAP_46_56);
			MULT_57(45)<=signed(DIN_57_7)*signed(FMAP_46_57);
			MULT_58(45)<=signed(DIN_58_7)*signed(FMAP_46_58);
			MULT_59(45)<=signed(DIN_59_7)*signed(FMAP_46_59);
			MULT_60(45)<=signed(DIN_60_7)*signed(FMAP_46_60);
			MULT_61(45)<=signed(DIN_61_7)*signed(FMAP_46_61);
			MULT_62(45)<=signed(DIN_62_7)*signed(FMAP_46_62);
			MULT_63(45)<=signed(DIN_63_7)*signed(FMAP_46_63);
			MULT_64(45)<=signed(DIN_64_7)*signed(FMAP_46_64);
			MULT_65(45)<=signed(DIN_65_7)*signed(FMAP_46_65);
			MULT_66(45)<=signed(DIN_66_7)*signed(FMAP_46_66);
			MULT_67(45)<=signed(DIN_67_7)*signed(FMAP_46_67);
			MULT_68(45)<=signed(DIN_68_7)*signed(FMAP_46_68);
			MULT_69(45)<=signed(DIN_69_7)*signed(FMAP_46_69);
			MULT_70(45)<=signed(DIN_70_7)*signed(FMAP_46_70);
			MULT_71(45)<=signed(DIN_71_7)*signed(FMAP_46_71);
			MULT_72(45)<=signed(DIN_72_7)*signed(FMAP_46_72);
			MULT_73(45)<=signed(DIN_73_7)*signed(FMAP_46_73);
			MULT_74(45)<=signed(DIN_74_7)*signed(FMAP_46_74);
			MULT_75(45)<=signed(DIN_75_7)*signed(FMAP_46_75);
			MULT_76(45)<=signed(DIN_76_7)*signed(FMAP_46_76);
			MULT_77(45)<=signed(DIN_77_7)*signed(FMAP_46_77);
			MULT_78(45)<=signed(DIN_78_7)*signed(FMAP_46_78);
			MULT_79(45)<=signed(DIN_79_7)*signed(FMAP_46_79);
			MULT_80(45)<=signed(DIN_80_7)*signed(FMAP_46_80);
			MULT_81(45)<=signed(DIN_81_7)*signed(FMAP_46_81);
			MULT_82(45)<=signed(DIN_82_7)*signed(FMAP_46_82);
			MULT_83(45)<=signed(DIN_83_7)*signed(FMAP_46_83);
			MULT_84(45)<=signed(DIN_84_7)*signed(FMAP_46_84);
			MULT_85(45)<=signed(DIN_85_7)*signed(FMAP_46_85);
			MULT_86(45)<=signed(DIN_86_7)*signed(FMAP_46_86);
			MULT_87(45)<=signed(DIN_87_7)*signed(FMAP_46_87);
			MULT_88(45)<=signed(DIN_88_7)*signed(FMAP_46_88);
			MULT_89(45)<=signed(DIN_89_7)*signed(FMAP_46_89);
			MULT_90(45)<=signed(DIN_90_7)*signed(FMAP_46_90);
			MULT_91(45)<=signed(DIN_91_7)*signed(FMAP_46_91);
			MULT_92(45)<=signed(DIN_92_7)*signed(FMAP_46_92);
			MULT_93(45)<=signed(DIN_93_7)*signed(FMAP_46_93);
			MULT_94(45)<=signed(DIN_94_7)*signed(FMAP_46_94);
			MULT_95(45)<=signed(DIN_95_7)*signed(FMAP_46_95);
			MULT_96(45)<=signed(DIN_96_7)*signed(FMAP_46_96);
			MULT_97(45)<=signed(DIN_97_7)*signed(FMAP_46_97);
			MULT_98(45)<=signed(DIN_98_7)*signed(FMAP_46_98);
			MULT_99(45)<=signed(DIN_99_7)*signed(FMAP_46_99);
			MULT_100(45)<=signed(DIN_100_7)*signed(FMAP_46_100);
			MULT_101(45)<=signed(DIN_101_7)*signed(FMAP_46_101);
			MULT_102(45)<=signed(DIN_102_7)*signed(FMAP_46_102);
			MULT_103(45)<=signed(DIN_103_7)*signed(FMAP_46_103);
			MULT_104(45)<=signed(DIN_104_7)*signed(FMAP_46_104);
			MULT_105(45)<=signed(DIN_105_7)*signed(FMAP_46_105);
			MULT_106(45)<=signed(DIN_106_7)*signed(FMAP_46_106);
			MULT_107(45)<=signed(DIN_107_7)*signed(FMAP_46_107);
			MULT_108(45)<=signed(DIN_108_7)*signed(FMAP_46_108);
			MULT_109(45)<=signed(DIN_109_7)*signed(FMAP_46_109);
			MULT_110(45)<=signed(DIN_110_7)*signed(FMAP_46_110);
			MULT_111(45)<=signed(DIN_111_7)*signed(FMAP_46_111);
			MULT_112(45)<=signed(DIN_112_7)*signed(FMAP_46_112);
			MULT_113(45)<=signed(DIN_113_7)*signed(FMAP_46_113);
			MULT_114(45)<=signed(DIN_114_7)*signed(FMAP_46_114);
			MULT_115(45)<=signed(DIN_115_7)*signed(FMAP_46_115);
			MULT_116(45)<=signed(DIN_116_7)*signed(FMAP_46_116);
			MULT_117(45)<=signed(DIN_117_7)*signed(FMAP_46_117);
			MULT_118(45)<=signed(DIN_118_7)*signed(FMAP_46_118);
			MULT_119(45)<=signed(DIN_119_7)*signed(FMAP_46_119);
			MULT_120(45)<=signed(DIN_120_7)*signed(FMAP_46_120);

			MULT_1(46)<=signed(DIN_1_7)*signed(FMAP_47_1);
			MULT_2(46)<=signed(DIN_2_7)*signed(FMAP_47_2);
			MULT_3(46)<=signed(DIN_3_7)*signed(FMAP_47_3);
			MULT_4(46)<=signed(DIN_4_7)*signed(FMAP_47_4);
			MULT_5(46)<=signed(DIN_5_7)*signed(FMAP_47_5);
			MULT_6(46)<=signed(DIN_6_7)*signed(FMAP_47_6);
			MULT_7(46)<=signed(DIN_7_7)*signed(FMAP_47_7);
			MULT_8(46)<=signed(DIN_8_7)*signed(FMAP_47_8);
			MULT_9(46)<=signed(DIN_9_7)*signed(FMAP_47_9);
			MULT_10(46)<=signed(DIN_10_7)*signed(FMAP_47_10);
			MULT_11(46)<=signed(DIN_11_7)*signed(FMAP_47_11);
			MULT_12(46)<=signed(DIN_12_7)*signed(FMAP_47_12);
			MULT_13(46)<=signed(DIN_13_7)*signed(FMAP_47_13);
			MULT_14(46)<=signed(DIN_14_7)*signed(FMAP_47_14);
			MULT_15(46)<=signed(DIN_15_7)*signed(FMAP_47_15);
			MULT_16(46)<=signed(DIN_16_7)*signed(FMAP_47_16);
			MULT_17(46)<=signed(DIN_17_7)*signed(FMAP_47_17);
			MULT_18(46)<=signed(DIN_18_7)*signed(FMAP_47_18);
			MULT_19(46)<=signed(DIN_19_7)*signed(FMAP_47_19);
			MULT_20(46)<=signed(DIN_20_7)*signed(FMAP_47_20);
			MULT_21(46)<=signed(DIN_21_7)*signed(FMAP_47_21);
			MULT_22(46)<=signed(DIN_22_7)*signed(FMAP_47_22);
			MULT_23(46)<=signed(DIN_23_7)*signed(FMAP_47_23);
			MULT_24(46)<=signed(DIN_24_7)*signed(FMAP_47_24);
			MULT_25(46)<=signed(DIN_25_7)*signed(FMAP_47_25);
			MULT_26(46)<=signed(DIN_26_7)*signed(FMAP_47_26);
			MULT_27(46)<=signed(DIN_27_7)*signed(FMAP_47_27);
			MULT_28(46)<=signed(DIN_28_7)*signed(FMAP_47_28);
			MULT_29(46)<=signed(DIN_29_7)*signed(FMAP_47_29);
			MULT_30(46)<=signed(DIN_30_7)*signed(FMAP_47_30);
			MULT_31(46)<=signed(DIN_31_7)*signed(FMAP_47_31);
			MULT_32(46)<=signed(DIN_32_7)*signed(FMAP_47_32);
			MULT_33(46)<=signed(DIN_33_7)*signed(FMAP_47_33);
			MULT_34(46)<=signed(DIN_34_7)*signed(FMAP_47_34);
			MULT_35(46)<=signed(DIN_35_7)*signed(FMAP_47_35);
			MULT_36(46)<=signed(DIN_36_7)*signed(FMAP_47_36);
			MULT_37(46)<=signed(DIN_37_7)*signed(FMAP_47_37);
			MULT_38(46)<=signed(DIN_38_7)*signed(FMAP_47_38);
			MULT_39(46)<=signed(DIN_39_7)*signed(FMAP_47_39);
			MULT_40(46)<=signed(DIN_40_7)*signed(FMAP_47_40);
			MULT_41(46)<=signed(DIN_41_7)*signed(FMAP_47_41);
			MULT_42(46)<=signed(DIN_42_7)*signed(FMAP_47_42);
			MULT_43(46)<=signed(DIN_43_7)*signed(FMAP_47_43);
			MULT_44(46)<=signed(DIN_44_7)*signed(FMAP_47_44);
			MULT_45(46)<=signed(DIN_45_7)*signed(FMAP_47_45);
			MULT_46(46)<=signed(DIN_46_7)*signed(FMAP_47_46);
			MULT_47(46)<=signed(DIN_47_7)*signed(FMAP_47_47);
			MULT_48(46)<=signed(DIN_48_7)*signed(FMAP_47_48);
			MULT_49(46)<=signed(DIN_49_7)*signed(FMAP_47_49);
			MULT_50(46)<=signed(DIN_50_7)*signed(FMAP_47_50);
			MULT_51(46)<=signed(DIN_51_7)*signed(FMAP_47_51);
			MULT_52(46)<=signed(DIN_52_7)*signed(FMAP_47_52);
			MULT_53(46)<=signed(DIN_53_7)*signed(FMAP_47_53);
			MULT_54(46)<=signed(DIN_54_7)*signed(FMAP_47_54);
			MULT_55(46)<=signed(DIN_55_7)*signed(FMAP_47_55);
			MULT_56(46)<=signed(DIN_56_7)*signed(FMAP_47_56);
			MULT_57(46)<=signed(DIN_57_7)*signed(FMAP_47_57);
			MULT_58(46)<=signed(DIN_58_7)*signed(FMAP_47_58);
			MULT_59(46)<=signed(DIN_59_7)*signed(FMAP_47_59);
			MULT_60(46)<=signed(DIN_60_7)*signed(FMAP_47_60);
			MULT_61(46)<=signed(DIN_61_7)*signed(FMAP_47_61);
			MULT_62(46)<=signed(DIN_62_7)*signed(FMAP_47_62);
			MULT_63(46)<=signed(DIN_63_7)*signed(FMAP_47_63);
			MULT_64(46)<=signed(DIN_64_7)*signed(FMAP_47_64);
			MULT_65(46)<=signed(DIN_65_7)*signed(FMAP_47_65);
			MULT_66(46)<=signed(DIN_66_7)*signed(FMAP_47_66);
			MULT_67(46)<=signed(DIN_67_7)*signed(FMAP_47_67);
			MULT_68(46)<=signed(DIN_68_7)*signed(FMAP_47_68);
			MULT_69(46)<=signed(DIN_69_7)*signed(FMAP_47_69);
			MULT_70(46)<=signed(DIN_70_7)*signed(FMAP_47_70);
			MULT_71(46)<=signed(DIN_71_7)*signed(FMAP_47_71);
			MULT_72(46)<=signed(DIN_72_7)*signed(FMAP_47_72);
			MULT_73(46)<=signed(DIN_73_7)*signed(FMAP_47_73);
			MULT_74(46)<=signed(DIN_74_7)*signed(FMAP_47_74);
			MULT_75(46)<=signed(DIN_75_7)*signed(FMAP_47_75);
			MULT_76(46)<=signed(DIN_76_7)*signed(FMAP_47_76);
			MULT_77(46)<=signed(DIN_77_7)*signed(FMAP_47_77);
			MULT_78(46)<=signed(DIN_78_7)*signed(FMAP_47_78);
			MULT_79(46)<=signed(DIN_79_7)*signed(FMAP_47_79);
			MULT_80(46)<=signed(DIN_80_7)*signed(FMAP_47_80);
			MULT_81(46)<=signed(DIN_81_7)*signed(FMAP_47_81);
			MULT_82(46)<=signed(DIN_82_7)*signed(FMAP_47_82);
			MULT_83(46)<=signed(DIN_83_7)*signed(FMAP_47_83);
			MULT_84(46)<=signed(DIN_84_7)*signed(FMAP_47_84);
			MULT_85(46)<=signed(DIN_85_7)*signed(FMAP_47_85);
			MULT_86(46)<=signed(DIN_86_7)*signed(FMAP_47_86);
			MULT_87(46)<=signed(DIN_87_7)*signed(FMAP_47_87);
			MULT_88(46)<=signed(DIN_88_7)*signed(FMAP_47_88);
			MULT_89(46)<=signed(DIN_89_7)*signed(FMAP_47_89);
			MULT_90(46)<=signed(DIN_90_7)*signed(FMAP_47_90);
			MULT_91(46)<=signed(DIN_91_7)*signed(FMAP_47_91);
			MULT_92(46)<=signed(DIN_92_7)*signed(FMAP_47_92);
			MULT_93(46)<=signed(DIN_93_7)*signed(FMAP_47_93);
			MULT_94(46)<=signed(DIN_94_7)*signed(FMAP_47_94);
			MULT_95(46)<=signed(DIN_95_7)*signed(FMAP_47_95);
			MULT_96(46)<=signed(DIN_96_7)*signed(FMAP_47_96);
			MULT_97(46)<=signed(DIN_97_7)*signed(FMAP_47_97);
			MULT_98(46)<=signed(DIN_98_7)*signed(FMAP_47_98);
			MULT_99(46)<=signed(DIN_99_7)*signed(FMAP_47_99);
			MULT_100(46)<=signed(DIN_100_7)*signed(FMAP_47_100);
			MULT_101(46)<=signed(DIN_101_7)*signed(FMAP_47_101);
			MULT_102(46)<=signed(DIN_102_7)*signed(FMAP_47_102);
			MULT_103(46)<=signed(DIN_103_7)*signed(FMAP_47_103);
			MULT_104(46)<=signed(DIN_104_7)*signed(FMAP_47_104);
			MULT_105(46)<=signed(DIN_105_7)*signed(FMAP_47_105);
			MULT_106(46)<=signed(DIN_106_7)*signed(FMAP_47_106);
			MULT_107(46)<=signed(DIN_107_7)*signed(FMAP_47_107);
			MULT_108(46)<=signed(DIN_108_7)*signed(FMAP_47_108);
			MULT_109(46)<=signed(DIN_109_7)*signed(FMAP_47_109);
			MULT_110(46)<=signed(DIN_110_7)*signed(FMAP_47_110);
			MULT_111(46)<=signed(DIN_111_7)*signed(FMAP_47_111);
			MULT_112(46)<=signed(DIN_112_7)*signed(FMAP_47_112);
			MULT_113(46)<=signed(DIN_113_7)*signed(FMAP_47_113);
			MULT_114(46)<=signed(DIN_114_7)*signed(FMAP_47_114);
			MULT_115(46)<=signed(DIN_115_7)*signed(FMAP_47_115);
			MULT_116(46)<=signed(DIN_116_7)*signed(FMAP_47_116);
			MULT_117(46)<=signed(DIN_117_7)*signed(FMAP_47_117);
			MULT_118(46)<=signed(DIN_118_7)*signed(FMAP_47_118);
			MULT_119(46)<=signed(DIN_119_7)*signed(FMAP_47_119);
			MULT_120(46)<=signed(DIN_120_7)*signed(FMAP_47_120);

			MULT_1(47)<=signed(DIN_1_7)*signed(FMAP_48_1);
			MULT_2(47)<=signed(DIN_2_7)*signed(FMAP_48_2);
			MULT_3(47)<=signed(DIN_3_7)*signed(FMAP_48_3);
			MULT_4(47)<=signed(DIN_4_7)*signed(FMAP_48_4);
			MULT_5(47)<=signed(DIN_5_7)*signed(FMAP_48_5);
			MULT_6(47)<=signed(DIN_6_7)*signed(FMAP_48_6);
			MULT_7(47)<=signed(DIN_7_7)*signed(FMAP_48_7);
			MULT_8(47)<=signed(DIN_8_7)*signed(FMAP_48_8);
			MULT_9(47)<=signed(DIN_9_7)*signed(FMAP_48_9);
			MULT_10(47)<=signed(DIN_10_7)*signed(FMAP_48_10);
			MULT_11(47)<=signed(DIN_11_7)*signed(FMAP_48_11);
			MULT_12(47)<=signed(DIN_12_7)*signed(FMAP_48_12);
			MULT_13(47)<=signed(DIN_13_7)*signed(FMAP_48_13);
			MULT_14(47)<=signed(DIN_14_7)*signed(FMAP_48_14);
			MULT_15(47)<=signed(DIN_15_7)*signed(FMAP_48_15);
			MULT_16(47)<=signed(DIN_16_7)*signed(FMAP_48_16);
			MULT_17(47)<=signed(DIN_17_7)*signed(FMAP_48_17);
			MULT_18(47)<=signed(DIN_18_7)*signed(FMAP_48_18);
			MULT_19(47)<=signed(DIN_19_7)*signed(FMAP_48_19);
			MULT_20(47)<=signed(DIN_20_7)*signed(FMAP_48_20);
			MULT_21(47)<=signed(DIN_21_7)*signed(FMAP_48_21);
			MULT_22(47)<=signed(DIN_22_7)*signed(FMAP_48_22);
			MULT_23(47)<=signed(DIN_23_7)*signed(FMAP_48_23);
			MULT_24(47)<=signed(DIN_24_7)*signed(FMAP_48_24);
			MULT_25(47)<=signed(DIN_25_7)*signed(FMAP_48_25);
			MULT_26(47)<=signed(DIN_26_7)*signed(FMAP_48_26);
			MULT_27(47)<=signed(DIN_27_7)*signed(FMAP_48_27);
			MULT_28(47)<=signed(DIN_28_7)*signed(FMAP_48_28);
			MULT_29(47)<=signed(DIN_29_7)*signed(FMAP_48_29);
			MULT_30(47)<=signed(DIN_30_7)*signed(FMAP_48_30);
			MULT_31(47)<=signed(DIN_31_7)*signed(FMAP_48_31);
			MULT_32(47)<=signed(DIN_32_7)*signed(FMAP_48_32);
			MULT_33(47)<=signed(DIN_33_7)*signed(FMAP_48_33);
			MULT_34(47)<=signed(DIN_34_7)*signed(FMAP_48_34);
			MULT_35(47)<=signed(DIN_35_7)*signed(FMAP_48_35);
			MULT_36(47)<=signed(DIN_36_7)*signed(FMAP_48_36);
			MULT_37(47)<=signed(DIN_37_7)*signed(FMAP_48_37);
			MULT_38(47)<=signed(DIN_38_7)*signed(FMAP_48_38);
			MULT_39(47)<=signed(DIN_39_7)*signed(FMAP_48_39);
			MULT_40(47)<=signed(DIN_40_7)*signed(FMAP_48_40);
			MULT_41(47)<=signed(DIN_41_7)*signed(FMAP_48_41);
			MULT_42(47)<=signed(DIN_42_7)*signed(FMAP_48_42);
			MULT_43(47)<=signed(DIN_43_7)*signed(FMAP_48_43);
			MULT_44(47)<=signed(DIN_44_7)*signed(FMAP_48_44);
			MULT_45(47)<=signed(DIN_45_7)*signed(FMAP_48_45);
			MULT_46(47)<=signed(DIN_46_7)*signed(FMAP_48_46);
			MULT_47(47)<=signed(DIN_47_7)*signed(FMAP_48_47);
			MULT_48(47)<=signed(DIN_48_7)*signed(FMAP_48_48);
			MULT_49(47)<=signed(DIN_49_7)*signed(FMAP_48_49);
			MULT_50(47)<=signed(DIN_50_7)*signed(FMAP_48_50);
			MULT_51(47)<=signed(DIN_51_7)*signed(FMAP_48_51);
			MULT_52(47)<=signed(DIN_52_7)*signed(FMAP_48_52);
			MULT_53(47)<=signed(DIN_53_7)*signed(FMAP_48_53);
			MULT_54(47)<=signed(DIN_54_7)*signed(FMAP_48_54);
			MULT_55(47)<=signed(DIN_55_7)*signed(FMAP_48_55);
			MULT_56(47)<=signed(DIN_56_7)*signed(FMAP_48_56);
			MULT_57(47)<=signed(DIN_57_7)*signed(FMAP_48_57);
			MULT_58(47)<=signed(DIN_58_7)*signed(FMAP_48_58);
			MULT_59(47)<=signed(DIN_59_7)*signed(FMAP_48_59);
			MULT_60(47)<=signed(DIN_60_7)*signed(FMAP_48_60);
			MULT_61(47)<=signed(DIN_61_7)*signed(FMAP_48_61);
			MULT_62(47)<=signed(DIN_62_7)*signed(FMAP_48_62);
			MULT_63(47)<=signed(DIN_63_7)*signed(FMAP_48_63);
			MULT_64(47)<=signed(DIN_64_7)*signed(FMAP_48_64);
			MULT_65(47)<=signed(DIN_65_7)*signed(FMAP_48_65);
			MULT_66(47)<=signed(DIN_66_7)*signed(FMAP_48_66);
			MULT_67(47)<=signed(DIN_67_7)*signed(FMAP_48_67);
			MULT_68(47)<=signed(DIN_68_7)*signed(FMAP_48_68);
			MULT_69(47)<=signed(DIN_69_7)*signed(FMAP_48_69);
			MULT_70(47)<=signed(DIN_70_7)*signed(FMAP_48_70);
			MULT_71(47)<=signed(DIN_71_7)*signed(FMAP_48_71);
			MULT_72(47)<=signed(DIN_72_7)*signed(FMAP_48_72);
			MULT_73(47)<=signed(DIN_73_7)*signed(FMAP_48_73);
			MULT_74(47)<=signed(DIN_74_7)*signed(FMAP_48_74);
			MULT_75(47)<=signed(DIN_75_7)*signed(FMAP_48_75);
			MULT_76(47)<=signed(DIN_76_7)*signed(FMAP_48_76);
			MULT_77(47)<=signed(DIN_77_7)*signed(FMAP_48_77);
			MULT_78(47)<=signed(DIN_78_7)*signed(FMAP_48_78);
			MULT_79(47)<=signed(DIN_79_7)*signed(FMAP_48_79);
			MULT_80(47)<=signed(DIN_80_7)*signed(FMAP_48_80);
			MULT_81(47)<=signed(DIN_81_7)*signed(FMAP_48_81);
			MULT_82(47)<=signed(DIN_82_7)*signed(FMAP_48_82);
			MULT_83(47)<=signed(DIN_83_7)*signed(FMAP_48_83);
			MULT_84(47)<=signed(DIN_84_7)*signed(FMAP_48_84);
			MULT_85(47)<=signed(DIN_85_7)*signed(FMAP_48_85);
			MULT_86(47)<=signed(DIN_86_7)*signed(FMAP_48_86);
			MULT_87(47)<=signed(DIN_87_7)*signed(FMAP_48_87);
			MULT_88(47)<=signed(DIN_88_7)*signed(FMAP_48_88);
			MULT_89(47)<=signed(DIN_89_7)*signed(FMAP_48_89);
			MULT_90(47)<=signed(DIN_90_7)*signed(FMAP_48_90);
			MULT_91(47)<=signed(DIN_91_7)*signed(FMAP_48_91);
			MULT_92(47)<=signed(DIN_92_7)*signed(FMAP_48_92);
			MULT_93(47)<=signed(DIN_93_7)*signed(FMAP_48_93);
			MULT_94(47)<=signed(DIN_94_7)*signed(FMAP_48_94);
			MULT_95(47)<=signed(DIN_95_7)*signed(FMAP_48_95);
			MULT_96(47)<=signed(DIN_96_7)*signed(FMAP_48_96);
			MULT_97(47)<=signed(DIN_97_7)*signed(FMAP_48_97);
			MULT_98(47)<=signed(DIN_98_7)*signed(FMAP_48_98);
			MULT_99(47)<=signed(DIN_99_7)*signed(FMAP_48_99);
			MULT_100(47)<=signed(DIN_100_7)*signed(FMAP_48_100);
			MULT_101(47)<=signed(DIN_101_7)*signed(FMAP_48_101);
			MULT_102(47)<=signed(DIN_102_7)*signed(FMAP_48_102);
			MULT_103(47)<=signed(DIN_103_7)*signed(FMAP_48_103);
			MULT_104(47)<=signed(DIN_104_7)*signed(FMAP_48_104);
			MULT_105(47)<=signed(DIN_105_7)*signed(FMAP_48_105);
			MULT_106(47)<=signed(DIN_106_7)*signed(FMAP_48_106);
			MULT_107(47)<=signed(DIN_107_7)*signed(FMAP_48_107);
			MULT_108(47)<=signed(DIN_108_7)*signed(FMAP_48_108);
			MULT_109(47)<=signed(DIN_109_7)*signed(FMAP_48_109);
			MULT_110(47)<=signed(DIN_110_7)*signed(FMAP_48_110);
			MULT_111(47)<=signed(DIN_111_7)*signed(FMAP_48_111);
			MULT_112(47)<=signed(DIN_112_7)*signed(FMAP_48_112);
			MULT_113(47)<=signed(DIN_113_7)*signed(FMAP_48_113);
			MULT_114(47)<=signed(DIN_114_7)*signed(FMAP_48_114);
			MULT_115(47)<=signed(DIN_115_7)*signed(FMAP_48_115);
			MULT_116(47)<=signed(DIN_116_7)*signed(FMAP_48_116);
			MULT_117(47)<=signed(DIN_117_7)*signed(FMAP_48_117);
			MULT_118(47)<=signed(DIN_118_7)*signed(FMAP_48_118);
			MULT_119(47)<=signed(DIN_119_7)*signed(FMAP_48_119);
			MULT_120(47)<=signed(DIN_120_7)*signed(FMAP_48_120);

			MULT_1(48)<=signed(DIN_1_7)*signed(FMAP_49_1);
			MULT_2(48)<=signed(DIN_2_7)*signed(FMAP_49_2);
			MULT_3(48)<=signed(DIN_3_7)*signed(FMAP_49_3);
			MULT_4(48)<=signed(DIN_4_7)*signed(FMAP_49_4);
			MULT_5(48)<=signed(DIN_5_7)*signed(FMAP_49_5);
			MULT_6(48)<=signed(DIN_6_7)*signed(FMAP_49_6);
			MULT_7(48)<=signed(DIN_7_7)*signed(FMAP_49_7);
			MULT_8(48)<=signed(DIN_8_7)*signed(FMAP_49_8);
			MULT_9(48)<=signed(DIN_9_7)*signed(FMAP_49_9);
			MULT_10(48)<=signed(DIN_10_7)*signed(FMAP_49_10);
			MULT_11(48)<=signed(DIN_11_7)*signed(FMAP_49_11);
			MULT_12(48)<=signed(DIN_12_7)*signed(FMAP_49_12);
			MULT_13(48)<=signed(DIN_13_7)*signed(FMAP_49_13);
			MULT_14(48)<=signed(DIN_14_7)*signed(FMAP_49_14);
			MULT_15(48)<=signed(DIN_15_7)*signed(FMAP_49_15);
			MULT_16(48)<=signed(DIN_16_7)*signed(FMAP_49_16);
			MULT_17(48)<=signed(DIN_17_7)*signed(FMAP_49_17);
			MULT_18(48)<=signed(DIN_18_7)*signed(FMAP_49_18);
			MULT_19(48)<=signed(DIN_19_7)*signed(FMAP_49_19);
			MULT_20(48)<=signed(DIN_20_7)*signed(FMAP_49_20);
			MULT_21(48)<=signed(DIN_21_7)*signed(FMAP_49_21);
			MULT_22(48)<=signed(DIN_22_7)*signed(FMAP_49_22);
			MULT_23(48)<=signed(DIN_23_7)*signed(FMAP_49_23);
			MULT_24(48)<=signed(DIN_24_7)*signed(FMAP_49_24);
			MULT_25(48)<=signed(DIN_25_7)*signed(FMAP_49_25);
			MULT_26(48)<=signed(DIN_26_7)*signed(FMAP_49_26);
			MULT_27(48)<=signed(DIN_27_7)*signed(FMAP_49_27);
			MULT_28(48)<=signed(DIN_28_7)*signed(FMAP_49_28);
			MULT_29(48)<=signed(DIN_29_7)*signed(FMAP_49_29);
			MULT_30(48)<=signed(DIN_30_7)*signed(FMAP_49_30);
			MULT_31(48)<=signed(DIN_31_7)*signed(FMAP_49_31);
			MULT_32(48)<=signed(DIN_32_7)*signed(FMAP_49_32);
			MULT_33(48)<=signed(DIN_33_7)*signed(FMAP_49_33);
			MULT_34(48)<=signed(DIN_34_7)*signed(FMAP_49_34);
			MULT_35(48)<=signed(DIN_35_7)*signed(FMAP_49_35);
			MULT_36(48)<=signed(DIN_36_7)*signed(FMAP_49_36);
			MULT_37(48)<=signed(DIN_37_7)*signed(FMAP_49_37);
			MULT_38(48)<=signed(DIN_38_7)*signed(FMAP_49_38);
			MULT_39(48)<=signed(DIN_39_7)*signed(FMAP_49_39);
			MULT_40(48)<=signed(DIN_40_7)*signed(FMAP_49_40);
			MULT_41(48)<=signed(DIN_41_7)*signed(FMAP_49_41);
			MULT_42(48)<=signed(DIN_42_7)*signed(FMAP_49_42);
			MULT_43(48)<=signed(DIN_43_7)*signed(FMAP_49_43);
			MULT_44(48)<=signed(DIN_44_7)*signed(FMAP_49_44);
			MULT_45(48)<=signed(DIN_45_7)*signed(FMAP_49_45);
			MULT_46(48)<=signed(DIN_46_7)*signed(FMAP_49_46);
			MULT_47(48)<=signed(DIN_47_7)*signed(FMAP_49_47);
			MULT_48(48)<=signed(DIN_48_7)*signed(FMAP_49_48);
			MULT_49(48)<=signed(DIN_49_7)*signed(FMAP_49_49);
			MULT_50(48)<=signed(DIN_50_7)*signed(FMAP_49_50);
			MULT_51(48)<=signed(DIN_51_7)*signed(FMAP_49_51);
			MULT_52(48)<=signed(DIN_52_7)*signed(FMAP_49_52);
			MULT_53(48)<=signed(DIN_53_7)*signed(FMAP_49_53);
			MULT_54(48)<=signed(DIN_54_7)*signed(FMAP_49_54);
			MULT_55(48)<=signed(DIN_55_7)*signed(FMAP_49_55);
			MULT_56(48)<=signed(DIN_56_7)*signed(FMAP_49_56);
			MULT_57(48)<=signed(DIN_57_7)*signed(FMAP_49_57);
			MULT_58(48)<=signed(DIN_58_7)*signed(FMAP_49_58);
			MULT_59(48)<=signed(DIN_59_7)*signed(FMAP_49_59);
			MULT_60(48)<=signed(DIN_60_7)*signed(FMAP_49_60);
			MULT_61(48)<=signed(DIN_61_7)*signed(FMAP_49_61);
			MULT_62(48)<=signed(DIN_62_7)*signed(FMAP_49_62);
			MULT_63(48)<=signed(DIN_63_7)*signed(FMAP_49_63);
			MULT_64(48)<=signed(DIN_64_7)*signed(FMAP_49_64);
			MULT_65(48)<=signed(DIN_65_7)*signed(FMAP_49_65);
			MULT_66(48)<=signed(DIN_66_7)*signed(FMAP_49_66);
			MULT_67(48)<=signed(DIN_67_7)*signed(FMAP_49_67);
			MULT_68(48)<=signed(DIN_68_7)*signed(FMAP_49_68);
			MULT_69(48)<=signed(DIN_69_7)*signed(FMAP_49_69);
			MULT_70(48)<=signed(DIN_70_7)*signed(FMAP_49_70);
			MULT_71(48)<=signed(DIN_71_7)*signed(FMAP_49_71);
			MULT_72(48)<=signed(DIN_72_7)*signed(FMAP_49_72);
			MULT_73(48)<=signed(DIN_73_7)*signed(FMAP_49_73);
			MULT_74(48)<=signed(DIN_74_7)*signed(FMAP_49_74);
			MULT_75(48)<=signed(DIN_75_7)*signed(FMAP_49_75);
			MULT_76(48)<=signed(DIN_76_7)*signed(FMAP_49_76);
			MULT_77(48)<=signed(DIN_77_7)*signed(FMAP_49_77);
			MULT_78(48)<=signed(DIN_78_7)*signed(FMAP_49_78);
			MULT_79(48)<=signed(DIN_79_7)*signed(FMAP_49_79);
			MULT_80(48)<=signed(DIN_80_7)*signed(FMAP_49_80);
			MULT_81(48)<=signed(DIN_81_7)*signed(FMAP_49_81);
			MULT_82(48)<=signed(DIN_82_7)*signed(FMAP_49_82);
			MULT_83(48)<=signed(DIN_83_7)*signed(FMAP_49_83);
			MULT_84(48)<=signed(DIN_84_7)*signed(FMAP_49_84);
			MULT_85(48)<=signed(DIN_85_7)*signed(FMAP_49_85);
			MULT_86(48)<=signed(DIN_86_7)*signed(FMAP_49_86);
			MULT_87(48)<=signed(DIN_87_7)*signed(FMAP_49_87);
			MULT_88(48)<=signed(DIN_88_7)*signed(FMAP_49_88);
			MULT_89(48)<=signed(DIN_89_7)*signed(FMAP_49_89);
			MULT_90(48)<=signed(DIN_90_7)*signed(FMAP_49_90);
			MULT_91(48)<=signed(DIN_91_7)*signed(FMAP_49_91);
			MULT_92(48)<=signed(DIN_92_7)*signed(FMAP_49_92);
			MULT_93(48)<=signed(DIN_93_7)*signed(FMAP_49_93);
			MULT_94(48)<=signed(DIN_94_7)*signed(FMAP_49_94);
			MULT_95(48)<=signed(DIN_95_7)*signed(FMAP_49_95);
			MULT_96(48)<=signed(DIN_96_7)*signed(FMAP_49_96);
			MULT_97(48)<=signed(DIN_97_7)*signed(FMAP_49_97);
			MULT_98(48)<=signed(DIN_98_7)*signed(FMAP_49_98);
			MULT_99(48)<=signed(DIN_99_7)*signed(FMAP_49_99);
			MULT_100(48)<=signed(DIN_100_7)*signed(FMAP_49_100);
			MULT_101(48)<=signed(DIN_101_7)*signed(FMAP_49_101);
			MULT_102(48)<=signed(DIN_102_7)*signed(FMAP_49_102);
			MULT_103(48)<=signed(DIN_103_7)*signed(FMAP_49_103);
			MULT_104(48)<=signed(DIN_104_7)*signed(FMAP_49_104);
			MULT_105(48)<=signed(DIN_105_7)*signed(FMAP_49_105);
			MULT_106(48)<=signed(DIN_106_7)*signed(FMAP_49_106);
			MULT_107(48)<=signed(DIN_107_7)*signed(FMAP_49_107);
			MULT_108(48)<=signed(DIN_108_7)*signed(FMAP_49_108);
			MULT_109(48)<=signed(DIN_109_7)*signed(FMAP_49_109);
			MULT_110(48)<=signed(DIN_110_7)*signed(FMAP_49_110);
			MULT_111(48)<=signed(DIN_111_7)*signed(FMAP_49_111);
			MULT_112(48)<=signed(DIN_112_7)*signed(FMAP_49_112);
			MULT_113(48)<=signed(DIN_113_7)*signed(FMAP_49_113);
			MULT_114(48)<=signed(DIN_114_7)*signed(FMAP_49_114);
			MULT_115(48)<=signed(DIN_115_7)*signed(FMAP_49_115);
			MULT_116(48)<=signed(DIN_116_7)*signed(FMAP_49_116);
			MULT_117(48)<=signed(DIN_117_7)*signed(FMAP_49_117);
			MULT_118(48)<=signed(DIN_118_7)*signed(FMAP_49_118);
			MULT_119(48)<=signed(DIN_119_7)*signed(FMAP_49_119);
			MULT_120(48)<=signed(DIN_120_7)*signed(FMAP_49_120);

			MULT_1(49)<=signed(DIN_1_7)*signed(FMAP_50_1);
			MULT_2(49)<=signed(DIN_2_7)*signed(FMAP_50_2);
			MULT_3(49)<=signed(DIN_3_7)*signed(FMAP_50_3);
			MULT_4(49)<=signed(DIN_4_7)*signed(FMAP_50_4);
			MULT_5(49)<=signed(DIN_5_7)*signed(FMAP_50_5);
			MULT_6(49)<=signed(DIN_6_7)*signed(FMAP_50_6);
			MULT_7(49)<=signed(DIN_7_7)*signed(FMAP_50_7);
			MULT_8(49)<=signed(DIN_8_7)*signed(FMAP_50_8);
			MULT_9(49)<=signed(DIN_9_7)*signed(FMAP_50_9);
			MULT_10(49)<=signed(DIN_10_7)*signed(FMAP_50_10);
			MULT_11(49)<=signed(DIN_11_7)*signed(FMAP_50_11);
			MULT_12(49)<=signed(DIN_12_7)*signed(FMAP_50_12);
			MULT_13(49)<=signed(DIN_13_7)*signed(FMAP_50_13);
			MULT_14(49)<=signed(DIN_14_7)*signed(FMAP_50_14);
			MULT_15(49)<=signed(DIN_15_7)*signed(FMAP_50_15);
			MULT_16(49)<=signed(DIN_16_7)*signed(FMAP_50_16);
			MULT_17(49)<=signed(DIN_17_7)*signed(FMAP_50_17);
			MULT_18(49)<=signed(DIN_18_7)*signed(FMAP_50_18);
			MULT_19(49)<=signed(DIN_19_7)*signed(FMAP_50_19);
			MULT_20(49)<=signed(DIN_20_7)*signed(FMAP_50_20);
			MULT_21(49)<=signed(DIN_21_7)*signed(FMAP_50_21);
			MULT_22(49)<=signed(DIN_22_7)*signed(FMAP_50_22);
			MULT_23(49)<=signed(DIN_23_7)*signed(FMAP_50_23);
			MULT_24(49)<=signed(DIN_24_7)*signed(FMAP_50_24);
			MULT_25(49)<=signed(DIN_25_7)*signed(FMAP_50_25);
			MULT_26(49)<=signed(DIN_26_7)*signed(FMAP_50_26);
			MULT_27(49)<=signed(DIN_27_7)*signed(FMAP_50_27);
			MULT_28(49)<=signed(DIN_28_7)*signed(FMAP_50_28);
			MULT_29(49)<=signed(DIN_29_7)*signed(FMAP_50_29);
			MULT_30(49)<=signed(DIN_30_7)*signed(FMAP_50_30);
			MULT_31(49)<=signed(DIN_31_7)*signed(FMAP_50_31);
			MULT_32(49)<=signed(DIN_32_7)*signed(FMAP_50_32);
			MULT_33(49)<=signed(DIN_33_7)*signed(FMAP_50_33);
			MULT_34(49)<=signed(DIN_34_7)*signed(FMAP_50_34);
			MULT_35(49)<=signed(DIN_35_7)*signed(FMAP_50_35);
			MULT_36(49)<=signed(DIN_36_7)*signed(FMAP_50_36);
			MULT_37(49)<=signed(DIN_37_7)*signed(FMAP_50_37);
			MULT_38(49)<=signed(DIN_38_7)*signed(FMAP_50_38);
			MULT_39(49)<=signed(DIN_39_7)*signed(FMAP_50_39);
			MULT_40(49)<=signed(DIN_40_7)*signed(FMAP_50_40);
			MULT_41(49)<=signed(DIN_41_7)*signed(FMAP_50_41);
			MULT_42(49)<=signed(DIN_42_7)*signed(FMAP_50_42);
			MULT_43(49)<=signed(DIN_43_7)*signed(FMAP_50_43);
			MULT_44(49)<=signed(DIN_44_7)*signed(FMAP_50_44);
			MULT_45(49)<=signed(DIN_45_7)*signed(FMAP_50_45);
			MULT_46(49)<=signed(DIN_46_7)*signed(FMAP_50_46);
			MULT_47(49)<=signed(DIN_47_7)*signed(FMAP_50_47);
			MULT_48(49)<=signed(DIN_48_7)*signed(FMAP_50_48);
			MULT_49(49)<=signed(DIN_49_7)*signed(FMAP_50_49);
			MULT_50(49)<=signed(DIN_50_7)*signed(FMAP_50_50);
			MULT_51(49)<=signed(DIN_51_7)*signed(FMAP_50_51);
			MULT_52(49)<=signed(DIN_52_7)*signed(FMAP_50_52);
			MULT_53(49)<=signed(DIN_53_7)*signed(FMAP_50_53);
			MULT_54(49)<=signed(DIN_54_7)*signed(FMAP_50_54);
			MULT_55(49)<=signed(DIN_55_7)*signed(FMAP_50_55);
			MULT_56(49)<=signed(DIN_56_7)*signed(FMAP_50_56);
			MULT_57(49)<=signed(DIN_57_7)*signed(FMAP_50_57);
			MULT_58(49)<=signed(DIN_58_7)*signed(FMAP_50_58);
			MULT_59(49)<=signed(DIN_59_7)*signed(FMAP_50_59);
			MULT_60(49)<=signed(DIN_60_7)*signed(FMAP_50_60);
			MULT_61(49)<=signed(DIN_61_7)*signed(FMAP_50_61);
			MULT_62(49)<=signed(DIN_62_7)*signed(FMAP_50_62);
			MULT_63(49)<=signed(DIN_63_7)*signed(FMAP_50_63);
			MULT_64(49)<=signed(DIN_64_7)*signed(FMAP_50_64);
			MULT_65(49)<=signed(DIN_65_7)*signed(FMAP_50_65);
			MULT_66(49)<=signed(DIN_66_7)*signed(FMAP_50_66);
			MULT_67(49)<=signed(DIN_67_7)*signed(FMAP_50_67);
			MULT_68(49)<=signed(DIN_68_7)*signed(FMAP_50_68);
			MULT_69(49)<=signed(DIN_69_7)*signed(FMAP_50_69);
			MULT_70(49)<=signed(DIN_70_7)*signed(FMAP_50_70);
			MULT_71(49)<=signed(DIN_71_7)*signed(FMAP_50_71);
			MULT_72(49)<=signed(DIN_72_7)*signed(FMAP_50_72);
			MULT_73(49)<=signed(DIN_73_7)*signed(FMAP_50_73);
			MULT_74(49)<=signed(DIN_74_7)*signed(FMAP_50_74);
			MULT_75(49)<=signed(DIN_75_7)*signed(FMAP_50_75);
			MULT_76(49)<=signed(DIN_76_7)*signed(FMAP_50_76);
			MULT_77(49)<=signed(DIN_77_7)*signed(FMAP_50_77);
			MULT_78(49)<=signed(DIN_78_7)*signed(FMAP_50_78);
			MULT_79(49)<=signed(DIN_79_7)*signed(FMAP_50_79);
			MULT_80(49)<=signed(DIN_80_7)*signed(FMAP_50_80);
			MULT_81(49)<=signed(DIN_81_7)*signed(FMAP_50_81);
			MULT_82(49)<=signed(DIN_82_7)*signed(FMAP_50_82);
			MULT_83(49)<=signed(DIN_83_7)*signed(FMAP_50_83);
			MULT_84(49)<=signed(DIN_84_7)*signed(FMAP_50_84);
			MULT_85(49)<=signed(DIN_85_7)*signed(FMAP_50_85);
			MULT_86(49)<=signed(DIN_86_7)*signed(FMAP_50_86);
			MULT_87(49)<=signed(DIN_87_7)*signed(FMAP_50_87);
			MULT_88(49)<=signed(DIN_88_7)*signed(FMAP_50_88);
			MULT_89(49)<=signed(DIN_89_7)*signed(FMAP_50_89);
			MULT_90(49)<=signed(DIN_90_7)*signed(FMAP_50_90);
			MULT_91(49)<=signed(DIN_91_7)*signed(FMAP_50_91);
			MULT_92(49)<=signed(DIN_92_7)*signed(FMAP_50_92);
			MULT_93(49)<=signed(DIN_93_7)*signed(FMAP_50_93);
			MULT_94(49)<=signed(DIN_94_7)*signed(FMAP_50_94);
			MULT_95(49)<=signed(DIN_95_7)*signed(FMAP_50_95);
			MULT_96(49)<=signed(DIN_96_7)*signed(FMAP_50_96);
			MULT_97(49)<=signed(DIN_97_7)*signed(FMAP_50_97);
			MULT_98(49)<=signed(DIN_98_7)*signed(FMAP_50_98);
			MULT_99(49)<=signed(DIN_99_7)*signed(FMAP_50_99);
			MULT_100(49)<=signed(DIN_100_7)*signed(FMAP_50_100);
			MULT_101(49)<=signed(DIN_101_7)*signed(FMAP_50_101);
			MULT_102(49)<=signed(DIN_102_7)*signed(FMAP_50_102);
			MULT_103(49)<=signed(DIN_103_7)*signed(FMAP_50_103);
			MULT_104(49)<=signed(DIN_104_7)*signed(FMAP_50_104);
			MULT_105(49)<=signed(DIN_105_7)*signed(FMAP_50_105);
			MULT_106(49)<=signed(DIN_106_7)*signed(FMAP_50_106);
			MULT_107(49)<=signed(DIN_107_7)*signed(FMAP_50_107);
			MULT_108(49)<=signed(DIN_108_7)*signed(FMAP_50_108);
			MULT_109(49)<=signed(DIN_109_7)*signed(FMAP_50_109);
			MULT_110(49)<=signed(DIN_110_7)*signed(FMAP_50_110);
			MULT_111(49)<=signed(DIN_111_7)*signed(FMAP_50_111);
			MULT_112(49)<=signed(DIN_112_7)*signed(FMAP_50_112);
			MULT_113(49)<=signed(DIN_113_7)*signed(FMAP_50_113);
			MULT_114(49)<=signed(DIN_114_7)*signed(FMAP_50_114);
			MULT_115(49)<=signed(DIN_115_7)*signed(FMAP_50_115);
			MULT_116(49)<=signed(DIN_116_7)*signed(FMAP_50_116);
			MULT_117(49)<=signed(DIN_117_7)*signed(FMAP_50_117);
			MULT_118(49)<=signed(DIN_118_7)*signed(FMAP_50_118);
			MULT_119(49)<=signed(DIN_119_7)*signed(FMAP_50_119);
			MULT_120(49)<=signed(DIN_120_7)*signed(FMAP_50_120);

			MULT_1(50)<=signed(DIN_1_7)*signed(FMAP_51_1);
			MULT_2(50)<=signed(DIN_2_7)*signed(FMAP_51_2);
			MULT_3(50)<=signed(DIN_3_7)*signed(FMAP_51_3);
			MULT_4(50)<=signed(DIN_4_7)*signed(FMAP_51_4);
			MULT_5(50)<=signed(DIN_5_7)*signed(FMAP_51_5);
			MULT_6(50)<=signed(DIN_6_7)*signed(FMAP_51_6);
			MULT_7(50)<=signed(DIN_7_7)*signed(FMAP_51_7);
			MULT_8(50)<=signed(DIN_8_7)*signed(FMAP_51_8);
			MULT_9(50)<=signed(DIN_9_7)*signed(FMAP_51_9);
			MULT_10(50)<=signed(DIN_10_7)*signed(FMAP_51_10);
			MULT_11(50)<=signed(DIN_11_7)*signed(FMAP_51_11);
			MULT_12(50)<=signed(DIN_12_7)*signed(FMAP_51_12);
			MULT_13(50)<=signed(DIN_13_7)*signed(FMAP_51_13);
			MULT_14(50)<=signed(DIN_14_7)*signed(FMAP_51_14);
			MULT_15(50)<=signed(DIN_15_7)*signed(FMAP_51_15);
			MULT_16(50)<=signed(DIN_16_7)*signed(FMAP_51_16);
			MULT_17(50)<=signed(DIN_17_7)*signed(FMAP_51_17);
			MULT_18(50)<=signed(DIN_18_7)*signed(FMAP_51_18);
			MULT_19(50)<=signed(DIN_19_7)*signed(FMAP_51_19);
			MULT_20(50)<=signed(DIN_20_7)*signed(FMAP_51_20);
			MULT_21(50)<=signed(DIN_21_7)*signed(FMAP_51_21);
			MULT_22(50)<=signed(DIN_22_7)*signed(FMAP_51_22);
			MULT_23(50)<=signed(DIN_23_7)*signed(FMAP_51_23);
			MULT_24(50)<=signed(DIN_24_7)*signed(FMAP_51_24);
			MULT_25(50)<=signed(DIN_25_7)*signed(FMAP_51_25);
			MULT_26(50)<=signed(DIN_26_7)*signed(FMAP_51_26);
			MULT_27(50)<=signed(DIN_27_7)*signed(FMAP_51_27);
			MULT_28(50)<=signed(DIN_28_7)*signed(FMAP_51_28);
			MULT_29(50)<=signed(DIN_29_7)*signed(FMAP_51_29);
			MULT_30(50)<=signed(DIN_30_7)*signed(FMAP_51_30);
			MULT_31(50)<=signed(DIN_31_7)*signed(FMAP_51_31);
			MULT_32(50)<=signed(DIN_32_7)*signed(FMAP_51_32);
			MULT_33(50)<=signed(DIN_33_7)*signed(FMAP_51_33);
			MULT_34(50)<=signed(DIN_34_7)*signed(FMAP_51_34);
			MULT_35(50)<=signed(DIN_35_7)*signed(FMAP_51_35);
			MULT_36(50)<=signed(DIN_36_7)*signed(FMAP_51_36);
			MULT_37(50)<=signed(DIN_37_7)*signed(FMAP_51_37);
			MULT_38(50)<=signed(DIN_38_7)*signed(FMAP_51_38);
			MULT_39(50)<=signed(DIN_39_7)*signed(FMAP_51_39);
			MULT_40(50)<=signed(DIN_40_7)*signed(FMAP_51_40);
			MULT_41(50)<=signed(DIN_41_7)*signed(FMAP_51_41);
			MULT_42(50)<=signed(DIN_42_7)*signed(FMAP_51_42);
			MULT_43(50)<=signed(DIN_43_7)*signed(FMAP_51_43);
			MULT_44(50)<=signed(DIN_44_7)*signed(FMAP_51_44);
			MULT_45(50)<=signed(DIN_45_7)*signed(FMAP_51_45);
			MULT_46(50)<=signed(DIN_46_7)*signed(FMAP_51_46);
			MULT_47(50)<=signed(DIN_47_7)*signed(FMAP_51_47);
			MULT_48(50)<=signed(DIN_48_7)*signed(FMAP_51_48);
			MULT_49(50)<=signed(DIN_49_7)*signed(FMAP_51_49);
			MULT_50(50)<=signed(DIN_50_7)*signed(FMAP_51_50);
			MULT_51(50)<=signed(DIN_51_7)*signed(FMAP_51_51);
			MULT_52(50)<=signed(DIN_52_7)*signed(FMAP_51_52);
			MULT_53(50)<=signed(DIN_53_7)*signed(FMAP_51_53);
			MULT_54(50)<=signed(DIN_54_7)*signed(FMAP_51_54);
			MULT_55(50)<=signed(DIN_55_7)*signed(FMAP_51_55);
			MULT_56(50)<=signed(DIN_56_7)*signed(FMAP_51_56);
			MULT_57(50)<=signed(DIN_57_7)*signed(FMAP_51_57);
			MULT_58(50)<=signed(DIN_58_7)*signed(FMAP_51_58);
			MULT_59(50)<=signed(DIN_59_7)*signed(FMAP_51_59);
			MULT_60(50)<=signed(DIN_60_7)*signed(FMAP_51_60);
			MULT_61(50)<=signed(DIN_61_7)*signed(FMAP_51_61);
			MULT_62(50)<=signed(DIN_62_7)*signed(FMAP_51_62);
			MULT_63(50)<=signed(DIN_63_7)*signed(FMAP_51_63);
			MULT_64(50)<=signed(DIN_64_7)*signed(FMAP_51_64);
			MULT_65(50)<=signed(DIN_65_7)*signed(FMAP_51_65);
			MULT_66(50)<=signed(DIN_66_7)*signed(FMAP_51_66);
			MULT_67(50)<=signed(DIN_67_7)*signed(FMAP_51_67);
			MULT_68(50)<=signed(DIN_68_7)*signed(FMAP_51_68);
			MULT_69(50)<=signed(DIN_69_7)*signed(FMAP_51_69);
			MULT_70(50)<=signed(DIN_70_7)*signed(FMAP_51_70);
			MULT_71(50)<=signed(DIN_71_7)*signed(FMAP_51_71);
			MULT_72(50)<=signed(DIN_72_7)*signed(FMAP_51_72);
			MULT_73(50)<=signed(DIN_73_7)*signed(FMAP_51_73);
			MULT_74(50)<=signed(DIN_74_7)*signed(FMAP_51_74);
			MULT_75(50)<=signed(DIN_75_7)*signed(FMAP_51_75);
			MULT_76(50)<=signed(DIN_76_7)*signed(FMAP_51_76);
			MULT_77(50)<=signed(DIN_77_7)*signed(FMAP_51_77);
			MULT_78(50)<=signed(DIN_78_7)*signed(FMAP_51_78);
			MULT_79(50)<=signed(DIN_79_7)*signed(FMAP_51_79);
			MULT_80(50)<=signed(DIN_80_7)*signed(FMAP_51_80);
			MULT_81(50)<=signed(DIN_81_7)*signed(FMAP_51_81);
			MULT_82(50)<=signed(DIN_82_7)*signed(FMAP_51_82);
			MULT_83(50)<=signed(DIN_83_7)*signed(FMAP_51_83);
			MULT_84(50)<=signed(DIN_84_7)*signed(FMAP_51_84);
			MULT_85(50)<=signed(DIN_85_7)*signed(FMAP_51_85);
			MULT_86(50)<=signed(DIN_86_7)*signed(FMAP_51_86);
			MULT_87(50)<=signed(DIN_87_7)*signed(FMAP_51_87);
			MULT_88(50)<=signed(DIN_88_7)*signed(FMAP_51_88);
			MULT_89(50)<=signed(DIN_89_7)*signed(FMAP_51_89);
			MULT_90(50)<=signed(DIN_90_7)*signed(FMAP_51_90);
			MULT_91(50)<=signed(DIN_91_7)*signed(FMAP_51_91);
			MULT_92(50)<=signed(DIN_92_7)*signed(FMAP_51_92);
			MULT_93(50)<=signed(DIN_93_7)*signed(FMAP_51_93);
			MULT_94(50)<=signed(DIN_94_7)*signed(FMAP_51_94);
			MULT_95(50)<=signed(DIN_95_7)*signed(FMAP_51_95);
			MULT_96(50)<=signed(DIN_96_7)*signed(FMAP_51_96);
			MULT_97(50)<=signed(DIN_97_7)*signed(FMAP_51_97);
			MULT_98(50)<=signed(DIN_98_7)*signed(FMAP_51_98);
			MULT_99(50)<=signed(DIN_99_7)*signed(FMAP_51_99);
			MULT_100(50)<=signed(DIN_100_7)*signed(FMAP_51_100);
			MULT_101(50)<=signed(DIN_101_7)*signed(FMAP_51_101);
			MULT_102(50)<=signed(DIN_102_7)*signed(FMAP_51_102);
			MULT_103(50)<=signed(DIN_103_7)*signed(FMAP_51_103);
			MULT_104(50)<=signed(DIN_104_7)*signed(FMAP_51_104);
			MULT_105(50)<=signed(DIN_105_7)*signed(FMAP_51_105);
			MULT_106(50)<=signed(DIN_106_7)*signed(FMAP_51_106);
			MULT_107(50)<=signed(DIN_107_7)*signed(FMAP_51_107);
			MULT_108(50)<=signed(DIN_108_7)*signed(FMAP_51_108);
			MULT_109(50)<=signed(DIN_109_7)*signed(FMAP_51_109);
			MULT_110(50)<=signed(DIN_110_7)*signed(FMAP_51_110);
			MULT_111(50)<=signed(DIN_111_7)*signed(FMAP_51_111);
			MULT_112(50)<=signed(DIN_112_7)*signed(FMAP_51_112);
			MULT_113(50)<=signed(DIN_113_7)*signed(FMAP_51_113);
			MULT_114(50)<=signed(DIN_114_7)*signed(FMAP_51_114);
			MULT_115(50)<=signed(DIN_115_7)*signed(FMAP_51_115);
			MULT_116(50)<=signed(DIN_116_7)*signed(FMAP_51_116);
			MULT_117(50)<=signed(DIN_117_7)*signed(FMAP_51_117);
			MULT_118(50)<=signed(DIN_118_7)*signed(FMAP_51_118);
			MULT_119(50)<=signed(DIN_119_7)*signed(FMAP_51_119);
			MULT_120(50)<=signed(DIN_120_7)*signed(FMAP_51_120);

			MULT_1(51)<=signed(DIN_1_7)*signed(FMAP_52_1);
			MULT_2(51)<=signed(DIN_2_7)*signed(FMAP_52_2);
			MULT_3(51)<=signed(DIN_3_7)*signed(FMAP_52_3);
			MULT_4(51)<=signed(DIN_4_7)*signed(FMAP_52_4);
			MULT_5(51)<=signed(DIN_5_7)*signed(FMAP_52_5);
			MULT_6(51)<=signed(DIN_6_7)*signed(FMAP_52_6);
			MULT_7(51)<=signed(DIN_7_7)*signed(FMAP_52_7);
			MULT_8(51)<=signed(DIN_8_7)*signed(FMAP_52_8);
			MULT_9(51)<=signed(DIN_9_7)*signed(FMAP_52_9);
			MULT_10(51)<=signed(DIN_10_7)*signed(FMAP_52_10);
			MULT_11(51)<=signed(DIN_11_7)*signed(FMAP_52_11);
			MULT_12(51)<=signed(DIN_12_7)*signed(FMAP_52_12);
			MULT_13(51)<=signed(DIN_13_7)*signed(FMAP_52_13);
			MULT_14(51)<=signed(DIN_14_7)*signed(FMAP_52_14);
			MULT_15(51)<=signed(DIN_15_7)*signed(FMAP_52_15);
			MULT_16(51)<=signed(DIN_16_7)*signed(FMAP_52_16);
			MULT_17(51)<=signed(DIN_17_7)*signed(FMAP_52_17);
			MULT_18(51)<=signed(DIN_18_7)*signed(FMAP_52_18);
			MULT_19(51)<=signed(DIN_19_7)*signed(FMAP_52_19);
			MULT_20(51)<=signed(DIN_20_7)*signed(FMAP_52_20);
			MULT_21(51)<=signed(DIN_21_7)*signed(FMAP_52_21);
			MULT_22(51)<=signed(DIN_22_7)*signed(FMAP_52_22);
			MULT_23(51)<=signed(DIN_23_7)*signed(FMAP_52_23);
			MULT_24(51)<=signed(DIN_24_7)*signed(FMAP_52_24);
			MULT_25(51)<=signed(DIN_25_7)*signed(FMAP_52_25);
			MULT_26(51)<=signed(DIN_26_7)*signed(FMAP_52_26);
			MULT_27(51)<=signed(DIN_27_7)*signed(FMAP_52_27);
			MULT_28(51)<=signed(DIN_28_7)*signed(FMAP_52_28);
			MULT_29(51)<=signed(DIN_29_7)*signed(FMAP_52_29);
			MULT_30(51)<=signed(DIN_30_7)*signed(FMAP_52_30);
			MULT_31(51)<=signed(DIN_31_7)*signed(FMAP_52_31);
			MULT_32(51)<=signed(DIN_32_7)*signed(FMAP_52_32);
			MULT_33(51)<=signed(DIN_33_7)*signed(FMAP_52_33);
			MULT_34(51)<=signed(DIN_34_7)*signed(FMAP_52_34);
			MULT_35(51)<=signed(DIN_35_7)*signed(FMAP_52_35);
			MULT_36(51)<=signed(DIN_36_7)*signed(FMAP_52_36);
			MULT_37(51)<=signed(DIN_37_7)*signed(FMAP_52_37);
			MULT_38(51)<=signed(DIN_38_7)*signed(FMAP_52_38);
			MULT_39(51)<=signed(DIN_39_7)*signed(FMAP_52_39);
			MULT_40(51)<=signed(DIN_40_7)*signed(FMAP_52_40);
			MULT_41(51)<=signed(DIN_41_7)*signed(FMAP_52_41);
			MULT_42(51)<=signed(DIN_42_7)*signed(FMAP_52_42);
			MULT_43(51)<=signed(DIN_43_7)*signed(FMAP_52_43);
			MULT_44(51)<=signed(DIN_44_7)*signed(FMAP_52_44);
			MULT_45(51)<=signed(DIN_45_7)*signed(FMAP_52_45);
			MULT_46(51)<=signed(DIN_46_7)*signed(FMAP_52_46);
			MULT_47(51)<=signed(DIN_47_7)*signed(FMAP_52_47);
			MULT_48(51)<=signed(DIN_48_7)*signed(FMAP_52_48);
			MULT_49(51)<=signed(DIN_49_7)*signed(FMAP_52_49);
			MULT_50(51)<=signed(DIN_50_7)*signed(FMAP_52_50);
			MULT_51(51)<=signed(DIN_51_7)*signed(FMAP_52_51);
			MULT_52(51)<=signed(DIN_52_7)*signed(FMAP_52_52);
			MULT_53(51)<=signed(DIN_53_7)*signed(FMAP_52_53);
			MULT_54(51)<=signed(DIN_54_7)*signed(FMAP_52_54);
			MULT_55(51)<=signed(DIN_55_7)*signed(FMAP_52_55);
			MULT_56(51)<=signed(DIN_56_7)*signed(FMAP_52_56);
			MULT_57(51)<=signed(DIN_57_7)*signed(FMAP_52_57);
			MULT_58(51)<=signed(DIN_58_7)*signed(FMAP_52_58);
			MULT_59(51)<=signed(DIN_59_7)*signed(FMAP_52_59);
			MULT_60(51)<=signed(DIN_60_7)*signed(FMAP_52_60);
			MULT_61(51)<=signed(DIN_61_7)*signed(FMAP_52_61);
			MULT_62(51)<=signed(DIN_62_7)*signed(FMAP_52_62);
			MULT_63(51)<=signed(DIN_63_7)*signed(FMAP_52_63);
			MULT_64(51)<=signed(DIN_64_7)*signed(FMAP_52_64);
			MULT_65(51)<=signed(DIN_65_7)*signed(FMAP_52_65);
			MULT_66(51)<=signed(DIN_66_7)*signed(FMAP_52_66);
			MULT_67(51)<=signed(DIN_67_7)*signed(FMAP_52_67);
			MULT_68(51)<=signed(DIN_68_7)*signed(FMAP_52_68);
			MULT_69(51)<=signed(DIN_69_7)*signed(FMAP_52_69);
			MULT_70(51)<=signed(DIN_70_7)*signed(FMAP_52_70);
			MULT_71(51)<=signed(DIN_71_7)*signed(FMAP_52_71);
			MULT_72(51)<=signed(DIN_72_7)*signed(FMAP_52_72);
			MULT_73(51)<=signed(DIN_73_7)*signed(FMAP_52_73);
			MULT_74(51)<=signed(DIN_74_7)*signed(FMAP_52_74);
			MULT_75(51)<=signed(DIN_75_7)*signed(FMAP_52_75);
			MULT_76(51)<=signed(DIN_76_7)*signed(FMAP_52_76);
			MULT_77(51)<=signed(DIN_77_7)*signed(FMAP_52_77);
			MULT_78(51)<=signed(DIN_78_7)*signed(FMAP_52_78);
			MULT_79(51)<=signed(DIN_79_7)*signed(FMAP_52_79);
			MULT_80(51)<=signed(DIN_80_7)*signed(FMAP_52_80);
			MULT_81(51)<=signed(DIN_81_7)*signed(FMAP_52_81);
			MULT_82(51)<=signed(DIN_82_7)*signed(FMAP_52_82);
			MULT_83(51)<=signed(DIN_83_7)*signed(FMAP_52_83);
			MULT_84(51)<=signed(DIN_84_7)*signed(FMAP_52_84);
			MULT_85(51)<=signed(DIN_85_7)*signed(FMAP_52_85);
			MULT_86(51)<=signed(DIN_86_7)*signed(FMAP_52_86);
			MULT_87(51)<=signed(DIN_87_7)*signed(FMAP_52_87);
			MULT_88(51)<=signed(DIN_88_7)*signed(FMAP_52_88);
			MULT_89(51)<=signed(DIN_89_7)*signed(FMAP_52_89);
			MULT_90(51)<=signed(DIN_90_7)*signed(FMAP_52_90);
			MULT_91(51)<=signed(DIN_91_7)*signed(FMAP_52_91);
			MULT_92(51)<=signed(DIN_92_7)*signed(FMAP_52_92);
			MULT_93(51)<=signed(DIN_93_7)*signed(FMAP_52_93);
			MULT_94(51)<=signed(DIN_94_7)*signed(FMAP_52_94);
			MULT_95(51)<=signed(DIN_95_7)*signed(FMAP_52_95);
			MULT_96(51)<=signed(DIN_96_7)*signed(FMAP_52_96);
			MULT_97(51)<=signed(DIN_97_7)*signed(FMAP_52_97);
			MULT_98(51)<=signed(DIN_98_7)*signed(FMAP_52_98);
			MULT_99(51)<=signed(DIN_99_7)*signed(FMAP_52_99);
			MULT_100(51)<=signed(DIN_100_7)*signed(FMAP_52_100);
			MULT_101(51)<=signed(DIN_101_7)*signed(FMAP_52_101);
			MULT_102(51)<=signed(DIN_102_7)*signed(FMAP_52_102);
			MULT_103(51)<=signed(DIN_103_7)*signed(FMAP_52_103);
			MULT_104(51)<=signed(DIN_104_7)*signed(FMAP_52_104);
			MULT_105(51)<=signed(DIN_105_7)*signed(FMAP_52_105);
			MULT_106(51)<=signed(DIN_106_7)*signed(FMAP_52_106);
			MULT_107(51)<=signed(DIN_107_7)*signed(FMAP_52_107);
			MULT_108(51)<=signed(DIN_108_7)*signed(FMAP_52_108);
			MULT_109(51)<=signed(DIN_109_7)*signed(FMAP_52_109);
			MULT_110(51)<=signed(DIN_110_7)*signed(FMAP_52_110);
			MULT_111(51)<=signed(DIN_111_7)*signed(FMAP_52_111);
			MULT_112(51)<=signed(DIN_112_7)*signed(FMAP_52_112);
			MULT_113(51)<=signed(DIN_113_7)*signed(FMAP_52_113);
			MULT_114(51)<=signed(DIN_114_7)*signed(FMAP_52_114);
			MULT_115(51)<=signed(DIN_115_7)*signed(FMAP_52_115);
			MULT_116(51)<=signed(DIN_116_7)*signed(FMAP_52_116);
			MULT_117(51)<=signed(DIN_117_7)*signed(FMAP_52_117);
			MULT_118(51)<=signed(DIN_118_7)*signed(FMAP_52_118);
			MULT_119(51)<=signed(DIN_119_7)*signed(FMAP_52_119);
			MULT_120(51)<=signed(DIN_120_7)*signed(FMAP_52_120);

			MULT_1(52)<=signed(DIN_1_7)*signed(FMAP_53_1);
			MULT_2(52)<=signed(DIN_2_7)*signed(FMAP_53_2);
			MULT_3(52)<=signed(DIN_3_7)*signed(FMAP_53_3);
			MULT_4(52)<=signed(DIN_4_7)*signed(FMAP_53_4);
			MULT_5(52)<=signed(DIN_5_7)*signed(FMAP_53_5);
			MULT_6(52)<=signed(DIN_6_7)*signed(FMAP_53_6);
			MULT_7(52)<=signed(DIN_7_7)*signed(FMAP_53_7);
			MULT_8(52)<=signed(DIN_8_7)*signed(FMAP_53_8);
			MULT_9(52)<=signed(DIN_9_7)*signed(FMAP_53_9);
			MULT_10(52)<=signed(DIN_10_7)*signed(FMAP_53_10);
			MULT_11(52)<=signed(DIN_11_7)*signed(FMAP_53_11);
			MULT_12(52)<=signed(DIN_12_7)*signed(FMAP_53_12);
			MULT_13(52)<=signed(DIN_13_7)*signed(FMAP_53_13);
			MULT_14(52)<=signed(DIN_14_7)*signed(FMAP_53_14);
			MULT_15(52)<=signed(DIN_15_7)*signed(FMAP_53_15);
			MULT_16(52)<=signed(DIN_16_7)*signed(FMAP_53_16);
			MULT_17(52)<=signed(DIN_17_7)*signed(FMAP_53_17);
			MULT_18(52)<=signed(DIN_18_7)*signed(FMAP_53_18);
			MULT_19(52)<=signed(DIN_19_7)*signed(FMAP_53_19);
			MULT_20(52)<=signed(DIN_20_7)*signed(FMAP_53_20);
			MULT_21(52)<=signed(DIN_21_7)*signed(FMAP_53_21);
			MULT_22(52)<=signed(DIN_22_7)*signed(FMAP_53_22);
			MULT_23(52)<=signed(DIN_23_7)*signed(FMAP_53_23);
			MULT_24(52)<=signed(DIN_24_7)*signed(FMAP_53_24);
			MULT_25(52)<=signed(DIN_25_7)*signed(FMAP_53_25);
			MULT_26(52)<=signed(DIN_26_7)*signed(FMAP_53_26);
			MULT_27(52)<=signed(DIN_27_7)*signed(FMAP_53_27);
			MULT_28(52)<=signed(DIN_28_7)*signed(FMAP_53_28);
			MULT_29(52)<=signed(DIN_29_7)*signed(FMAP_53_29);
			MULT_30(52)<=signed(DIN_30_7)*signed(FMAP_53_30);
			MULT_31(52)<=signed(DIN_31_7)*signed(FMAP_53_31);
			MULT_32(52)<=signed(DIN_32_7)*signed(FMAP_53_32);
			MULT_33(52)<=signed(DIN_33_7)*signed(FMAP_53_33);
			MULT_34(52)<=signed(DIN_34_7)*signed(FMAP_53_34);
			MULT_35(52)<=signed(DIN_35_7)*signed(FMAP_53_35);
			MULT_36(52)<=signed(DIN_36_7)*signed(FMAP_53_36);
			MULT_37(52)<=signed(DIN_37_7)*signed(FMAP_53_37);
			MULT_38(52)<=signed(DIN_38_7)*signed(FMAP_53_38);
			MULT_39(52)<=signed(DIN_39_7)*signed(FMAP_53_39);
			MULT_40(52)<=signed(DIN_40_7)*signed(FMAP_53_40);
			MULT_41(52)<=signed(DIN_41_7)*signed(FMAP_53_41);
			MULT_42(52)<=signed(DIN_42_7)*signed(FMAP_53_42);
			MULT_43(52)<=signed(DIN_43_7)*signed(FMAP_53_43);
			MULT_44(52)<=signed(DIN_44_7)*signed(FMAP_53_44);
			MULT_45(52)<=signed(DIN_45_7)*signed(FMAP_53_45);
			MULT_46(52)<=signed(DIN_46_7)*signed(FMAP_53_46);
			MULT_47(52)<=signed(DIN_47_7)*signed(FMAP_53_47);
			MULT_48(52)<=signed(DIN_48_7)*signed(FMAP_53_48);
			MULT_49(52)<=signed(DIN_49_7)*signed(FMAP_53_49);
			MULT_50(52)<=signed(DIN_50_7)*signed(FMAP_53_50);
			MULT_51(52)<=signed(DIN_51_7)*signed(FMAP_53_51);
			MULT_52(52)<=signed(DIN_52_7)*signed(FMAP_53_52);
			MULT_53(52)<=signed(DIN_53_7)*signed(FMAP_53_53);
			MULT_54(52)<=signed(DIN_54_7)*signed(FMAP_53_54);
			MULT_55(52)<=signed(DIN_55_7)*signed(FMAP_53_55);
			MULT_56(52)<=signed(DIN_56_7)*signed(FMAP_53_56);
			MULT_57(52)<=signed(DIN_57_7)*signed(FMAP_53_57);
			MULT_58(52)<=signed(DIN_58_7)*signed(FMAP_53_58);
			MULT_59(52)<=signed(DIN_59_7)*signed(FMAP_53_59);
			MULT_60(52)<=signed(DIN_60_7)*signed(FMAP_53_60);
			MULT_61(52)<=signed(DIN_61_7)*signed(FMAP_53_61);
			MULT_62(52)<=signed(DIN_62_7)*signed(FMAP_53_62);
			MULT_63(52)<=signed(DIN_63_7)*signed(FMAP_53_63);
			MULT_64(52)<=signed(DIN_64_7)*signed(FMAP_53_64);
			MULT_65(52)<=signed(DIN_65_7)*signed(FMAP_53_65);
			MULT_66(52)<=signed(DIN_66_7)*signed(FMAP_53_66);
			MULT_67(52)<=signed(DIN_67_7)*signed(FMAP_53_67);
			MULT_68(52)<=signed(DIN_68_7)*signed(FMAP_53_68);
			MULT_69(52)<=signed(DIN_69_7)*signed(FMAP_53_69);
			MULT_70(52)<=signed(DIN_70_7)*signed(FMAP_53_70);
			MULT_71(52)<=signed(DIN_71_7)*signed(FMAP_53_71);
			MULT_72(52)<=signed(DIN_72_7)*signed(FMAP_53_72);
			MULT_73(52)<=signed(DIN_73_7)*signed(FMAP_53_73);
			MULT_74(52)<=signed(DIN_74_7)*signed(FMAP_53_74);
			MULT_75(52)<=signed(DIN_75_7)*signed(FMAP_53_75);
			MULT_76(52)<=signed(DIN_76_7)*signed(FMAP_53_76);
			MULT_77(52)<=signed(DIN_77_7)*signed(FMAP_53_77);
			MULT_78(52)<=signed(DIN_78_7)*signed(FMAP_53_78);
			MULT_79(52)<=signed(DIN_79_7)*signed(FMAP_53_79);
			MULT_80(52)<=signed(DIN_80_7)*signed(FMAP_53_80);
			MULT_81(52)<=signed(DIN_81_7)*signed(FMAP_53_81);
			MULT_82(52)<=signed(DIN_82_7)*signed(FMAP_53_82);
			MULT_83(52)<=signed(DIN_83_7)*signed(FMAP_53_83);
			MULT_84(52)<=signed(DIN_84_7)*signed(FMAP_53_84);
			MULT_85(52)<=signed(DIN_85_7)*signed(FMAP_53_85);
			MULT_86(52)<=signed(DIN_86_7)*signed(FMAP_53_86);
			MULT_87(52)<=signed(DIN_87_7)*signed(FMAP_53_87);
			MULT_88(52)<=signed(DIN_88_7)*signed(FMAP_53_88);
			MULT_89(52)<=signed(DIN_89_7)*signed(FMAP_53_89);
			MULT_90(52)<=signed(DIN_90_7)*signed(FMAP_53_90);
			MULT_91(52)<=signed(DIN_91_7)*signed(FMAP_53_91);
			MULT_92(52)<=signed(DIN_92_7)*signed(FMAP_53_92);
			MULT_93(52)<=signed(DIN_93_7)*signed(FMAP_53_93);
			MULT_94(52)<=signed(DIN_94_7)*signed(FMAP_53_94);
			MULT_95(52)<=signed(DIN_95_7)*signed(FMAP_53_95);
			MULT_96(52)<=signed(DIN_96_7)*signed(FMAP_53_96);
			MULT_97(52)<=signed(DIN_97_7)*signed(FMAP_53_97);
			MULT_98(52)<=signed(DIN_98_7)*signed(FMAP_53_98);
			MULT_99(52)<=signed(DIN_99_7)*signed(FMAP_53_99);
			MULT_100(52)<=signed(DIN_100_7)*signed(FMAP_53_100);
			MULT_101(52)<=signed(DIN_101_7)*signed(FMAP_53_101);
			MULT_102(52)<=signed(DIN_102_7)*signed(FMAP_53_102);
			MULT_103(52)<=signed(DIN_103_7)*signed(FMAP_53_103);
			MULT_104(52)<=signed(DIN_104_7)*signed(FMAP_53_104);
			MULT_105(52)<=signed(DIN_105_7)*signed(FMAP_53_105);
			MULT_106(52)<=signed(DIN_106_7)*signed(FMAP_53_106);
			MULT_107(52)<=signed(DIN_107_7)*signed(FMAP_53_107);
			MULT_108(52)<=signed(DIN_108_7)*signed(FMAP_53_108);
			MULT_109(52)<=signed(DIN_109_7)*signed(FMAP_53_109);
			MULT_110(52)<=signed(DIN_110_7)*signed(FMAP_53_110);
			MULT_111(52)<=signed(DIN_111_7)*signed(FMAP_53_111);
			MULT_112(52)<=signed(DIN_112_7)*signed(FMAP_53_112);
			MULT_113(52)<=signed(DIN_113_7)*signed(FMAP_53_113);
			MULT_114(52)<=signed(DIN_114_7)*signed(FMAP_53_114);
			MULT_115(52)<=signed(DIN_115_7)*signed(FMAP_53_115);
			MULT_116(52)<=signed(DIN_116_7)*signed(FMAP_53_116);
			MULT_117(52)<=signed(DIN_117_7)*signed(FMAP_53_117);
			MULT_118(52)<=signed(DIN_118_7)*signed(FMAP_53_118);
			MULT_119(52)<=signed(DIN_119_7)*signed(FMAP_53_119);
			MULT_120(52)<=signed(DIN_120_7)*signed(FMAP_53_120);

			MULT_1(53)<=signed(DIN_1_7)*signed(FMAP_54_1);
			MULT_2(53)<=signed(DIN_2_7)*signed(FMAP_54_2);
			MULT_3(53)<=signed(DIN_3_7)*signed(FMAP_54_3);
			MULT_4(53)<=signed(DIN_4_7)*signed(FMAP_54_4);
			MULT_5(53)<=signed(DIN_5_7)*signed(FMAP_54_5);
			MULT_6(53)<=signed(DIN_6_7)*signed(FMAP_54_6);
			MULT_7(53)<=signed(DIN_7_7)*signed(FMAP_54_7);
			MULT_8(53)<=signed(DIN_8_7)*signed(FMAP_54_8);
			MULT_9(53)<=signed(DIN_9_7)*signed(FMAP_54_9);
			MULT_10(53)<=signed(DIN_10_7)*signed(FMAP_54_10);
			MULT_11(53)<=signed(DIN_11_7)*signed(FMAP_54_11);
			MULT_12(53)<=signed(DIN_12_7)*signed(FMAP_54_12);
			MULT_13(53)<=signed(DIN_13_7)*signed(FMAP_54_13);
			MULT_14(53)<=signed(DIN_14_7)*signed(FMAP_54_14);
			MULT_15(53)<=signed(DIN_15_7)*signed(FMAP_54_15);
			MULT_16(53)<=signed(DIN_16_7)*signed(FMAP_54_16);
			MULT_17(53)<=signed(DIN_17_7)*signed(FMAP_54_17);
			MULT_18(53)<=signed(DIN_18_7)*signed(FMAP_54_18);
			MULT_19(53)<=signed(DIN_19_7)*signed(FMAP_54_19);
			MULT_20(53)<=signed(DIN_20_7)*signed(FMAP_54_20);
			MULT_21(53)<=signed(DIN_21_7)*signed(FMAP_54_21);
			MULT_22(53)<=signed(DIN_22_7)*signed(FMAP_54_22);
			MULT_23(53)<=signed(DIN_23_7)*signed(FMAP_54_23);
			MULT_24(53)<=signed(DIN_24_7)*signed(FMAP_54_24);
			MULT_25(53)<=signed(DIN_25_7)*signed(FMAP_54_25);
			MULT_26(53)<=signed(DIN_26_7)*signed(FMAP_54_26);
			MULT_27(53)<=signed(DIN_27_7)*signed(FMAP_54_27);
			MULT_28(53)<=signed(DIN_28_7)*signed(FMAP_54_28);
			MULT_29(53)<=signed(DIN_29_7)*signed(FMAP_54_29);
			MULT_30(53)<=signed(DIN_30_7)*signed(FMAP_54_30);
			MULT_31(53)<=signed(DIN_31_7)*signed(FMAP_54_31);
			MULT_32(53)<=signed(DIN_32_7)*signed(FMAP_54_32);
			MULT_33(53)<=signed(DIN_33_7)*signed(FMAP_54_33);
			MULT_34(53)<=signed(DIN_34_7)*signed(FMAP_54_34);
			MULT_35(53)<=signed(DIN_35_7)*signed(FMAP_54_35);
			MULT_36(53)<=signed(DIN_36_7)*signed(FMAP_54_36);
			MULT_37(53)<=signed(DIN_37_7)*signed(FMAP_54_37);
			MULT_38(53)<=signed(DIN_38_7)*signed(FMAP_54_38);
			MULT_39(53)<=signed(DIN_39_7)*signed(FMAP_54_39);
			MULT_40(53)<=signed(DIN_40_7)*signed(FMAP_54_40);
			MULT_41(53)<=signed(DIN_41_7)*signed(FMAP_54_41);
			MULT_42(53)<=signed(DIN_42_7)*signed(FMAP_54_42);
			MULT_43(53)<=signed(DIN_43_7)*signed(FMAP_54_43);
			MULT_44(53)<=signed(DIN_44_7)*signed(FMAP_54_44);
			MULT_45(53)<=signed(DIN_45_7)*signed(FMAP_54_45);
			MULT_46(53)<=signed(DIN_46_7)*signed(FMAP_54_46);
			MULT_47(53)<=signed(DIN_47_7)*signed(FMAP_54_47);
			MULT_48(53)<=signed(DIN_48_7)*signed(FMAP_54_48);
			MULT_49(53)<=signed(DIN_49_7)*signed(FMAP_54_49);
			MULT_50(53)<=signed(DIN_50_7)*signed(FMAP_54_50);
			MULT_51(53)<=signed(DIN_51_7)*signed(FMAP_54_51);
			MULT_52(53)<=signed(DIN_52_7)*signed(FMAP_54_52);
			MULT_53(53)<=signed(DIN_53_7)*signed(FMAP_54_53);
			MULT_54(53)<=signed(DIN_54_7)*signed(FMAP_54_54);
			MULT_55(53)<=signed(DIN_55_7)*signed(FMAP_54_55);
			MULT_56(53)<=signed(DIN_56_7)*signed(FMAP_54_56);
			MULT_57(53)<=signed(DIN_57_7)*signed(FMAP_54_57);
			MULT_58(53)<=signed(DIN_58_7)*signed(FMAP_54_58);
			MULT_59(53)<=signed(DIN_59_7)*signed(FMAP_54_59);
			MULT_60(53)<=signed(DIN_60_7)*signed(FMAP_54_60);
			MULT_61(53)<=signed(DIN_61_7)*signed(FMAP_54_61);
			MULT_62(53)<=signed(DIN_62_7)*signed(FMAP_54_62);
			MULT_63(53)<=signed(DIN_63_7)*signed(FMAP_54_63);
			MULT_64(53)<=signed(DIN_64_7)*signed(FMAP_54_64);
			MULT_65(53)<=signed(DIN_65_7)*signed(FMAP_54_65);
			MULT_66(53)<=signed(DIN_66_7)*signed(FMAP_54_66);
			MULT_67(53)<=signed(DIN_67_7)*signed(FMAP_54_67);
			MULT_68(53)<=signed(DIN_68_7)*signed(FMAP_54_68);
			MULT_69(53)<=signed(DIN_69_7)*signed(FMAP_54_69);
			MULT_70(53)<=signed(DIN_70_7)*signed(FMAP_54_70);
			MULT_71(53)<=signed(DIN_71_7)*signed(FMAP_54_71);
			MULT_72(53)<=signed(DIN_72_7)*signed(FMAP_54_72);
			MULT_73(53)<=signed(DIN_73_7)*signed(FMAP_54_73);
			MULT_74(53)<=signed(DIN_74_7)*signed(FMAP_54_74);
			MULT_75(53)<=signed(DIN_75_7)*signed(FMAP_54_75);
			MULT_76(53)<=signed(DIN_76_7)*signed(FMAP_54_76);
			MULT_77(53)<=signed(DIN_77_7)*signed(FMAP_54_77);
			MULT_78(53)<=signed(DIN_78_7)*signed(FMAP_54_78);
			MULT_79(53)<=signed(DIN_79_7)*signed(FMAP_54_79);
			MULT_80(53)<=signed(DIN_80_7)*signed(FMAP_54_80);
			MULT_81(53)<=signed(DIN_81_7)*signed(FMAP_54_81);
			MULT_82(53)<=signed(DIN_82_7)*signed(FMAP_54_82);
			MULT_83(53)<=signed(DIN_83_7)*signed(FMAP_54_83);
			MULT_84(53)<=signed(DIN_84_7)*signed(FMAP_54_84);
			MULT_85(53)<=signed(DIN_85_7)*signed(FMAP_54_85);
			MULT_86(53)<=signed(DIN_86_7)*signed(FMAP_54_86);
			MULT_87(53)<=signed(DIN_87_7)*signed(FMAP_54_87);
			MULT_88(53)<=signed(DIN_88_7)*signed(FMAP_54_88);
			MULT_89(53)<=signed(DIN_89_7)*signed(FMAP_54_89);
			MULT_90(53)<=signed(DIN_90_7)*signed(FMAP_54_90);
			MULT_91(53)<=signed(DIN_91_7)*signed(FMAP_54_91);
			MULT_92(53)<=signed(DIN_92_7)*signed(FMAP_54_92);
			MULT_93(53)<=signed(DIN_93_7)*signed(FMAP_54_93);
			MULT_94(53)<=signed(DIN_94_7)*signed(FMAP_54_94);
			MULT_95(53)<=signed(DIN_95_7)*signed(FMAP_54_95);
			MULT_96(53)<=signed(DIN_96_7)*signed(FMAP_54_96);
			MULT_97(53)<=signed(DIN_97_7)*signed(FMAP_54_97);
			MULT_98(53)<=signed(DIN_98_7)*signed(FMAP_54_98);
			MULT_99(53)<=signed(DIN_99_7)*signed(FMAP_54_99);
			MULT_100(53)<=signed(DIN_100_7)*signed(FMAP_54_100);
			MULT_101(53)<=signed(DIN_101_7)*signed(FMAP_54_101);
			MULT_102(53)<=signed(DIN_102_7)*signed(FMAP_54_102);
			MULT_103(53)<=signed(DIN_103_7)*signed(FMAP_54_103);
			MULT_104(53)<=signed(DIN_104_7)*signed(FMAP_54_104);
			MULT_105(53)<=signed(DIN_105_7)*signed(FMAP_54_105);
			MULT_106(53)<=signed(DIN_106_7)*signed(FMAP_54_106);
			MULT_107(53)<=signed(DIN_107_7)*signed(FMAP_54_107);
			MULT_108(53)<=signed(DIN_108_7)*signed(FMAP_54_108);
			MULT_109(53)<=signed(DIN_109_7)*signed(FMAP_54_109);
			MULT_110(53)<=signed(DIN_110_7)*signed(FMAP_54_110);
			MULT_111(53)<=signed(DIN_111_7)*signed(FMAP_54_111);
			MULT_112(53)<=signed(DIN_112_7)*signed(FMAP_54_112);
			MULT_113(53)<=signed(DIN_113_7)*signed(FMAP_54_113);
			MULT_114(53)<=signed(DIN_114_7)*signed(FMAP_54_114);
			MULT_115(53)<=signed(DIN_115_7)*signed(FMAP_54_115);
			MULT_116(53)<=signed(DIN_116_7)*signed(FMAP_54_116);
			MULT_117(53)<=signed(DIN_117_7)*signed(FMAP_54_117);
			MULT_118(53)<=signed(DIN_118_7)*signed(FMAP_54_118);
			MULT_119(53)<=signed(DIN_119_7)*signed(FMAP_54_119);
			MULT_120(53)<=signed(DIN_120_7)*signed(FMAP_54_120);

			MULT_1(54)<=signed(DIN_1_7)*signed(FMAP_55_1);
			MULT_2(54)<=signed(DIN_2_7)*signed(FMAP_55_2);
			MULT_3(54)<=signed(DIN_3_7)*signed(FMAP_55_3);
			MULT_4(54)<=signed(DIN_4_7)*signed(FMAP_55_4);
			MULT_5(54)<=signed(DIN_5_7)*signed(FMAP_55_5);
			MULT_6(54)<=signed(DIN_6_7)*signed(FMAP_55_6);
			MULT_7(54)<=signed(DIN_7_7)*signed(FMAP_55_7);
			MULT_8(54)<=signed(DIN_8_7)*signed(FMAP_55_8);
			MULT_9(54)<=signed(DIN_9_7)*signed(FMAP_55_9);
			MULT_10(54)<=signed(DIN_10_7)*signed(FMAP_55_10);
			MULT_11(54)<=signed(DIN_11_7)*signed(FMAP_55_11);
			MULT_12(54)<=signed(DIN_12_7)*signed(FMAP_55_12);
			MULT_13(54)<=signed(DIN_13_7)*signed(FMAP_55_13);
			MULT_14(54)<=signed(DIN_14_7)*signed(FMAP_55_14);
			MULT_15(54)<=signed(DIN_15_7)*signed(FMAP_55_15);
			MULT_16(54)<=signed(DIN_16_7)*signed(FMAP_55_16);
			MULT_17(54)<=signed(DIN_17_7)*signed(FMAP_55_17);
			MULT_18(54)<=signed(DIN_18_7)*signed(FMAP_55_18);
			MULT_19(54)<=signed(DIN_19_7)*signed(FMAP_55_19);
			MULT_20(54)<=signed(DIN_20_7)*signed(FMAP_55_20);
			MULT_21(54)<=signed(DIN_21_7)*signed(FMAP_55_21);
			MULT_22(54)<=signed(DIN_22_7)*signed(FMAP_55_22);
			MULT_23(54)<=signed(DIN_23_7)*signed(FMAP_55_23);
			MULT_24(54)<=signed(DIN_24_7)*signed(FMAP_55_24);
			MULT_25(54)<=signed(DIN_25_7)*signed(FMAP_55_25);
			MULT_26(54)<=signed(DIN_26_7)*signed(FMAP_55_26);
			MULT_27(54)<=signed(DIN_27_7)*signed(FMAP_55_27);
			MULT_28(54)<=signed(DIN_28_7)*signed(FMAP_55_28);
			MULT_29(54)<=signed(DIN_29_7)*signed(FMAP_55_29);
			MULT_30(54)<=signed(DIN_30_7)*signed(FMAP_55_30);
			MULT_31(54)<=signed(DIN_31_7)*signed(FMAP_55_31);
			MULT_32(54)<=signed(DIN_32_7)*signed(FMAP_55_32);
			MULT_33(54)<=signed(DIN_33_7)*signed(FMAP_55_33);
			MULT_34(54)<=signed(DIN_34_7)*signed(FMAP_55_34);
			MULT_35(54)<=signed(DIN_35_7)*signed(FMAP_55_35);
			MULT_36(54)<=signed(DIN_36_7)*signed(FMAP_55_36);
			MULT_37(54)<=signed(DIN_37_7)*signed(FMAP_55_37);
			MULT_38(54)<=signed(DIN_38_7)*signed(FMAP_55_38);
			MULT_39(54)<=signed(DIN_39_7)*signed(FMAP_55_39);
			MULT_40(54)<=signed(DIN_40_7)*signed(FMAP_55_40);
			MULT_41(54)<=signed(DIN_41_7)*signed(FMAP_55_41);
			MULT_42(54)<=signed(DIN_42_7)*signed(FMAP_55_42);
			MULT_43(54)<=signed(DIN_43_7)*signed(FMAP_55_43);
			MULT_44(54)<=signed(DIN_44_7)*signed(FMAP_55_44);
			MULT_45(54)<=signed(DIN_45_7)*signed(FMAP_55_45);
			MULT_46(54)<=signed(DIN_46_7)*signed(FMAP_55_46);
			MULT_47(54)<=signed(DIN_47_7)*signed(FMAP_55_47);
			MULT_48(54)<=signed(DIN_48_7)*signed(FMAP_55_48);
			MULT_49(54)<=signed(DIN_49_7)*signed(FMAP_55_49);
			MULT_50(54)<=signed(DIN_50_7)*signed(FMAP_55_50);
			MULT_51(54)<=signed(DIN_51_7)*signed(FMAP_55_51);
			MULT_52(54)<=signed(DIN_52_7)*signed(FMAP_55_52);
			MULT_53(54)<=signed(DIN_53_7)*signed(FMAP_55_53);
			MULT_54(54)<=signed(DIN_54_7)*signed(FMAP_55_54);
			MULT_55(54)<=signed(DIN_55_7)*signed(FMAP_55_55);
			MULT_56(54)<=signed(DIN_56_7)*signed(FMAP_55_56);
			MULT_57(54)<=signed(DIN_57_7)*signed(FMAP_55_57);
			MULT_58(54)<=signed(DIN_58_7)*signed(FMAP_55_58);
			MULT_59(54)<=signed(DIN_59_7)*signed(FMAP_55_59);
			MULT_60(54)<=signed(DIN_60_7)*signed(FMAP_55_60);
			MULT_61(54)<=signed(DIN_61_7)*signed(FMAP_55_61);
			MULT_62(54)<=signed(DIN_62_7)*signed(FMAP_55_62);
			MULT_63(54)<=signed(DIN_63_7)*signed(FMAP_55_63);
			MULT_64(54)<=signed(DIN_64_7)*signed(FMAP_55_64);
			MULT_65(54)<=signed(DIN_65_7)*signed(FMAP_55_65);
			MULT_66(54)<=signed(DIN_66_7)*signed(FMAP_55_66);
			MULT_67(54)<=signed(DIN_67_7)*signed(FMAP_55_67);
			MULT_68(54)<=signed(DIN_68_7)*signed(FMAP_55_68);
			MULT_69(54)<=signed(DIN_69_7)*signed(FMAP_55_69);
			MULT_70(54)<=signed(DIN_70_7)*signed(FMAP_55_70);
			MULT_71(54)<=signed(DIN_71_7)*signed(FMAP_55_71);
			MULT_72(54)<=signed(DIN_72_7)*signed(FMAP_55_72);
			MULT_73(54)<=signed(DIN_73_7)*signed(FMAP_55_73);
			MULT_74(54)<=signed(DIN_74_7)*signed(FMAP_55_74);
			MULT_75(54)<=signed(DIN_75_7)*signed(FMAP_55_75);
			MULT_76(54)<=signed(DIN_76_7)*signed(FMAP_55_76);
			MULT_77(54)<=signed(DIN_77_7)*signed(FMAP_55_77);
			MULT_78(54)<=signed(DIN_78_7)*signed(FMAP_55_78);
			MULT_79(54)<=signed(DIN_79_7)*signed(FMAP_55_79);
			MULT_80(54)<=signed(DIN_80_7)*signed(FMAP_55_80);
			MULT_81(54)<=signed(DIN_81_7)*signed(FMAP_55_81);
			MULT_82(54)<=signed(DIN_82_7)*signed(FMAP_55_82);
			MULT_83(54)<=signed(DIN_83_7)*signed(FMAP_55_83);
			MULT_84(54)<=signed(DIN_84_7)*signed(FMAP_55_84);
			MULT_85(54)<=signed(DIN_85_7)*signed(FMAP_55_85);
			MULT_86(54)<=signed(DIN_86_7)*signed(FMAP_55_86);
			MULT_87(54)<=signed(DIN_87_7)*signed(FMAP_55_87);
			MULT_88(54)<=signed(DIN_88_7)*signed(FMAP_55_88);
			MULT_89(54)<=signed(DIN_89_7)*signed(FMAP_55_89);
			MULT_90(54)<=signed(DIN_90_7)*signed(FMAP_55_90);
			MULT_91(54)<=signed(DIN_91_7)*signed(FMAP_55_91);
			MULT_92(54)<=signed(DIN_92_7)*signed(FMAP_55_92);
			MULT_93(54)<=signed(DIN_93_7)*signed(FMAP_55_93);
			MULT_94(54)<=signed(DIN_94_7)*signed(FMAP_55_94);
			MULT_95(54)<=signed(DIN_95_7)*signed(FMAP_55_95);
			MULT_96(54)<=signed(DIN_96_7)*signed(FMAP_55_96);
			MULT_97(54)<=signed(DIN_97_7)*signed(FMAP_55_97);
			MULT_98(54)<=signed(DIN_98_7)*signed(FMAP_55_98);
			MULT_99(54)<=signed(DIN_99_7)*signed(FMAP_55_99);
			MULT_100(54)<=signed(DIN_100_7)*signed(FMAP_55_100);
			MULT_101(54)<=signed(DIN_101_7)*signed(FMAP_55_101);
			MULT_102(54)<=signed(DIN_102_7)*signed(FMAP_55_102);
			MULT_103(54)<=signed(DIN_103_7)*signed(FMAP_55_103);
			MULT_104(54)<=signed(DIN_104_7)*signed(FMAP_55_104);
			MULT_105(54)<=signed(DIN_105_7)*signed(FMAP_55_105);
			MULT_106(54)<=signed(DIN_106_7)*signed(FMAP_55_106);
			MULT_107(54)<=signed(DIN_107_7)*signed(FMAP_55_107);
			MULT_108(54)<=signed(DIN_108_7)*signed(FMAP_55_108);
			MULT_109(54)<=signed(DIN_109_7)*signed(FMAP_55_109);
			MULT_110(54)<=signed(DIN_110_7)*signed(FMAP_55_110);
			MULT_111(54)<=signed(DIN_111_7)*signed(FMAP_55_111);
			MULT_112(54)<=signed(DIN_112_7)*signed(FMAP_55_112);
			MULT_113(54)<=signed(DIN_113_7)*signed(FMAP_55_113);
			MULT_114(54)<=signed(DIN_114_7)*signed(FMAP_55_114);
			MULT_115(54)<=signed(DIN_115_7)*signed(FMAP_55_115);
			MULT_116(54)<=signed(DIN_116_7)*signed(FMAP_55_116);
			MULT_117(54)<=signed(DIN_117_7)*signed(FMAP_55_117);
			MULT_118(54)<=signed(DIN_118_7)*signed(FMAP_55_118);
			MULT_119(54)<=signed(DIN_119_7)*signed(FMAP_55_119);
			MULT_120(54)<=signed(DIN_120_7)*signed(FMAP_55_120);

			MULT_1(55)<=signed(DIN_1_7)*signed(FMAP_56_1);
			MULT_2(55)<=signed(DIN_2_7)*signed(FMAP_56_2);
			MULT_3(55)<=signed(DIN_3_7)*signed(FMAP_56_3);
			MULT_4(55)<=signed(DIN_4_7)*signed(FMAP_56_4);
			MULT_5(55)<=signed(DIN_5_7)*signed(FMAP_56_5);
			MULT_6(55)<=signed(DIN_6_7)*signed(FMAP_56_6);
			MULT_7(55)<=signed(DIN_7_7)*signed(FMAP_56_7);
			MULT_8(55)<=signed(DIN_8_7)*signed(FMAP_56_8);
			MULT_9(55)<=signed(DIN_9_7)*signed(FMAP_56_9);
			MULT_10(55)<=signed(DIN_10_7)*signed(FMAP_56_10);
			MULT_11(55)<=signed(DIN_11_7)*signed(FMAP_56_11);
			MULT_12(55)<=signed(DIN_12_7)*signed(FMAP_56_12);
			MULT_13(55)<=signed(DIN_13_7)*signed(FMAP_56_13);
			MULT_14(55)<=signed(DIN_14_7)*signed(FMAP_56_14);
			MULT_15(55)<=signed(DIN_15_7)*signed(FMAP_56_15);
			MULT_16(55)<=signed(DIN_16_7)*signed(FMAP_56_16);
			MULT_17(55)<=signed(DIN_17_7)*signed(FMAP_56_17);
			MULT_18(55)<=signed(DIN_18_7)*signed(FMAP_56_18);
			MULT_19(55)<=signed(DIN_19_7)*signed(FMAP_56_19);
			MULT_20(55)<=signed(DIN_20_7)*signed(FMAP_56_20);
			MULT_21(55)<=signed(DIN_21_7)*signed(FMAP_56_21);
			MULT_22(55)<=signed(DIN_22_7)*signed(FMAP_56_22);
			MULT_23(55)<=signed(DIN_23_7)*signed(FMAP_56_23);
			MULT_24(55)<=signed(DIN_24_7)*signed(FMAP_56_24);
			MULT_25(55)<=signed(DIN_25_7)*signed(FMAP_56_25);
			MULT_26(55)<=signed(DIN_26_7)*signed(FMAP_56_26);
			MULT_27(55)<=signed(DIN_27_7)*signed(FMAP_56_27);
			MULT_28(55)<=signed(DIN_28_7)*signed(FMAP_56_28);
			MULT_29(55)<=signed(DIN_29_7)*signed(FMAP_56_29);
			MULT_30(55)<=signed(DIN_30_7)*signed(FMAP_56_30);
			MULT_31(55)<=signed(DIN_31_7)*signed(FMAP_56_31);
			MULT_32(55)<=signed(DIN_32_7)*signed(FMAP_56_32);
			MULT_33(55)<=signed(DIN_33_7)*signed(FMAP_56_33);
			MULT_34(55)<=signed(DIN_34_7)*signed(FMAP_56_34);
			MULT_35(55)<=signed(DIN_35_7)*signed(FMAP_56_35);
			MULT_36(55)<=signed(DIN_36_7)*signed(FMAP_56_36);
			MULT_37(55)<=signed(DIN_37_7)*signed(FMAP_56_37);
			MULT_38(55)<=signed(DIN_38_7)*signed(FMAP_56_38);
			MULT_39(55)<=signed(DIN_39_7)*signed(FMAP_56_39);
			MULT_40(55)<=signed(DIN_40_7)*signed(FMAP_56_40);
			MULT_41(55)<=signed(DIN_41_7)*signed(FMAP_56_41);
			MULT_42(55)<=signed(DIN_42_7)*signed(FMAP_56_42);
			MULT_43(55)<=signed(DIN_43_7)*signed(FMAP_56_43);
			MULT_44(55)<=signed(DIN_44_7)*signed(FMAP_56_44);
			MULT_45(55)<=signed(DIN_45_7)*signed(FMAP_56_45);
			MULT_46(55)<=signed(DIN_46_7)*signed(FMAP_56_46);
			MULT_47(55)<=signed(DIN_47_7)*signed(FMAP_56_47);
			MULT_48(55)<=signed(DIN_48_7)*signed(FMAP_56_48);
			MULT_49(55)<=signed(DIN_49_7)*signed(FMAP_56_49);
			MULT_50(55)<=signed(DIN_50_7)*signed(FMAP_56_50);
			MULT_51(55)<=signed(DIN_51_7)*signed(FMAP_56_51);
			MULT_52(55)<=signed(DIN_52_7)*signed(FMAP_56_52);
			MULT_53(55)<=signed(DIN_53_7)*signed(FMAP_56_53);
			MULT_54(55)<=signed(DIN_54_7)*signed(FMAP_56_54);
			MULT_55(55)<=signed(DIN_55_7)*signed(FMAP_56_55);
			MULT_56(55)<=signed(DIN_56_7)*signed(FMAP_56_56);
			MULT_57(55)<=signed(DIN_57_7)*signed(FMAP_56_57);
			MULT_58(55)<=signed(DIN_58_7)*signed(FMAP_56_58);
			MULT_59(55)<=signed(DIN_59_7)*signed(FMAP_56_59);
			MULT_60(55)<=signed(DIN_60_7)*signed(FMAP_56_60);
			MULT_61(55)<=signed(DIN_61_7)*signed(FMAP_56_61);
			MULT_62(55)<=signed(DIN_62_7)*signed(FMAP_56_62);
			MULT_63(55)<=signed(DIN_63_7)*signed(FMAP_56_63);
			MULT_64(55)<=signed(DIN_64_7)*signed(FMAP_56_64);
			MULT_65(55)<=signed(DIN_65_7)*signed(FMAP_56_65);
			MULT_66(55)<=signed(DIN_66_7)*signed(FMAP_56_66);
			MULT_67(55)<=signed(DIN_67_7)*signed(FMAP_56_67);
			MULT_68(55)<=signed(DIN_68_7)*signed(FMAP_56_68);
			MULT_69(55)<=signed(DIN_69_7)*signed(FMAP_56_69);
			MULT_70(55)<=signed(DIN_70_7)*signed(FMAP_56_70);
			MULT_71(55)<=signed(DIN_71_7)*signed(FMAP_56_71);
			MULT_72(55)<=signed(DIN_72_7)*signed(FMAP_56_72);
			MULT_73(55)<=signed(DIN_73_7)*signed(FMAP_56_73);
			MULT_74(55)<=signed(DIN_74_7)*signed(FMAP_56_74);
			MULT_75(55)<=signed(DIN_75_7)*signed(FMAP_56_75);
			MULT_76(55)<=signed(DIN_76_7)*signed(FMAP_56_76);
			MULT_77(55)<=signed(DIN_77_7)*signed(FMAP_56_77);
			MULT_78(55)<=signed(DIN_78_7)*signed(FMAP_56_78);
			MULT_79(55)<=signed(DIN_79_7)*signed(FMAP_56_79);
			MULT_80(55)<=signed(DIN_80_7)*signed(FMAP_56_80);
			MULT_81(55)<=signed(DIN_81_7)*signed(FMAP_56_81);
			MULT_82(55)<=signed(DIN_82_7)*signed(FMAP_56_82);
			MULT_83(55)<=signed(DIN_83_7)*signed(FMAP_56_83);
			MULT_84(55)<=signed(DIN_84_7)*signed(FMAP_56_84);
			MULT_85(55)<=signed(DIN_85_7)*signed(FMAP_56_85);
			MULT_86(55)<=signed(DIN_86_7)*signed(FMAP_56_86);
			MULT_87(55)<=signed(DIN_87_7)*signed(FMAP_56_87);
			MULT_88(55)<=signed(DIN_88_7)*signed(FMAP_56_88);
			MULT_89(55)<=signed(DIN_89_7)*signed(FMAP_56_89);
			MULT_90(55)<=signed(DIN_90_7)*signed(FMAP_56_90);
			MULT_91(55)<=signed(DIN_91_7)*signed(FMAP_56_91);
			MULT_92(55)<=signed(DIN_92_7)*signed(FMAP_56_92);
			MULT_93(55)<=signed(DIN_93_7)*signed(FMAP_56_93);
			MULT_94(55)<=signed(DIN_94_7)*signed(FMAP_56_94);
			MULT_95(55)<=signed(DIN_95_7)*signed(FMAP_56_95);
			MULT_96(55)<=signed(DIN_96_7)*signed(FMAP_56_96);
			MULT_97(55)<=signed(DIN_97_7)*signed(FMAP_56_97);
			MULT_98(55)<=signed(DIN_98_7)*signed(FMAP_56_98);
			MULT_99(55)<=signed(DIN_99_7)*signed(FMAP_56_99);
			MULT_100(55)<=signed(DIN_100_7)*signed(FMAP_56_100);
			MULT_101(55)<=signed(DIN_101_7)*signed(FMAP_56_101);
			MULT_102(55)<=signed(DIN_102_7)*signed(FMAP_56_102);
			MULT_103(55)<=signed(DIN_103_7)*signed(FMAP_56_103);
			MULT_104(55)<=signed(DIN_104_7)*signed(FMAP_56_104);
			MULT_105(55)<=signed(DIN_105_7)*signed(FMAP_56_105);
			MULT_106(55)<=signed(DIN_106_7)*signed(FMAP_56_106);
			MULT_107(55)<=signed(DIN_107_7)*signed(FMAP_56_107);
			MULT_108(55)<=signed(DIN_108_7)*signed(FMAP_56_108);
			MULT_109(55)<=signed(DIN_109_7)*signed(FMAP_56_109);
			MULT_110(55)<=signed(DIN_110_7)*signed(FMAP_56_110);
			MULT_111(55)<=signed(DIN_111_7)*signed(FMAP_56_111);
			MULT_112(55)<=signed(DIN_112_7)*signed(FMAP_56_112);
			MULT_113(55)<=signed(DIN_113_7)*signed(FMAP_56_113);
			MULT_114(55)<=signed(DIN_114_7)*signed(FMAP_56_114);
			MULT_115(55)<=signed(DIN_115_7)*signed(FMAP_56_115);
			MULT_116(55)<=signed(DIN_116_7)*signed(FMAP_56_116);
			MULT_117(55)<=signed(DIN_117_7)*signed(FMAP_56_117);
			MULT_118(55)<=signed(DIN_118_7)*signed(FMAP_56_118);
			MULT_119(55)<=signed(DIN_119_7)*signed(FMAP_56_119);
			MULT_120(55)<=signed(DIN_120_7)*signed(FMAP_56_120);

			MULT_1(56)<=signed(DIN_1_7)*signed(FMAP_57_1);
			MULT_2(56)<=signed(DIN_2_7)*signed(FMAP_57_2);
			MULT_3(56)<=signed(DIN_3_7)*signed(FMAP_57_3);
			MULT_4(56)<=signed(DIN_4_7)*signed(FMAP_57_4);
			MULT_5(56)<=signed(DIN_5_7)*signed(FMAP_57_5);
			MULT_6(56)<=signed(DIN_6_7)*signed(FMAP_57_6);
			MULT_7(56)<=signed(DIN_7_7)*signed(FMAP_57_7);
			MULT_8(56)<=signed(DIN_8_7)*signed(FMAP_57_8);
			MULT_9(56)<=signed(DIN_9_7)*signed(FMAP_57_9);
			MULT_10(56)<=signed(DIN_10_7)*signed(FMAP_57_10);
			MULT_11(56)<=signed(DIN_11_7)*signed(FMAP_57_11);
			MULT_12(56)<=signed(DIN_12_7)*signed(FMAP_57_12);
			MULT_13(56)<=signed(DIN_13_7)*signed(FMAP_57_13);
			MULT_14(56)<=signed(DIN_14_7)*signed(FMAP_57_14);
			MULT_15(56)<=signed(DIN_15_7)*signed(FMAP_57_15);
			MULT_16(56)<=signed(DIN_16_7)*signed(FMAP_57_16);
			MULT_17(56)<=signed(DIN_17_7)*signed(FMAP_57_17);
			MULT_18(56)<=signed(DIN_18_7)*signed(FMAP_57_18);
			MULT_19(56)<=signed(DIN_19_7)*signed(FMAP_57_19);
			MULT_20(56)<=signed(DIN_20_7)*signed(FMAP_57_20);
			MULT_21(56)<=signed(DIN_21_7)*signed(FMAP_57_21);
			MULT_22(56)<=signed(DIN_22_7)*signed(FMAP_57_22);
			MULT_23(56)<=signed(DIN_23_7)*signed(FMAP_57_23);
			MULT_24(56)<=signed(DIN_24_7)*signed(FMAP_57_24);
			MULT_25(56)<=signed(DIN_25_7)*signed(FMAP_57_25);
			MULT_26(56)<=signed(DIN_26_7)*signed(FMAP_57_26);
			MULT_27(56)<=signed(DIN_27_7)*signed(FMAP_57_27);
			MULT_28(56)<=signed(DIN_28_7)*signed(FMAP_57_28);
			MULT_29(56)<=signed(DIN_29_7)*signed(FMAP_57_29);
			MULT_30(56)<=signed(DIN_30_7)*signed(FMAP_57_30);
			MULT_31(56)<=signed(DIN_31_7)*signed(FMAP_57_31);
			MULT_32(56)<=signed(DIN_32_7)*signed(FMAP_57_32);
			MULT_33(56)<=signed(DIN_33_7)*signed(FMAP_57_33);
			MULT_34(56)<=signed(DIN_34_7)*signed(FMAP_57_34);
			MULT_35(56)<=signed(DIN_35_7)*signed(FMAP_57_35);
			MULT_36(56)<=signed(DIN_36_7)*signed(FMAP_57_36);
			MULT_37(56)<=signed(DIN_37_7)*signed(FMAP_57_37);
			MULT_38(56)<=signed(DIN_38_7)*signed(FMAP_57_38);
			MULT_39(56)<=signed(DIN_39_7)*signed(FMAP_57_39);
			MULT_40(56)<=signed(DIN_40_7)*signed(FMAP_57_40);
			MULT_41(56)<=signed(DIN_41_7)*signed(FMAP_57_41);
			MULT_42(56)<=signed(DIN_42_7)*signed(FMAP_57_42);
			MULT_43(56)<=signed(DIN_43_7)*signed(FMAP_57_43);
			MULT_44(56)<=signed(DIN_44_7)*signed(FMAP_57_44);
			MULT_45(56)<=signed(DIN_45_7)*signed(FMAP_57_45);
			MULT_46(56)<=signed(DIN_46_7)*signed(FMAP_57_46);
			MULT_47(56)<=signed(DIN_47_7)*signed(FMAP_57_47);
			MULT_48(56)<=signed(DIN_48_7)*signed(FMAP_57_48);
			MULT_49(56)<=signed(DIN_49_7)*signed(FMAP_57_49);
			MULT_50(56)<=signed(DIN_50_7)*signed(FMAP_57_50);
			MULT_51(56)<=signed(DIN_51_7)*signed(FMAP_57_51);
			MULT_52(56)<=signed(DIN_52_7)*signed(FMAP_57_52);
			MULT_53(56)<=signed(DIN_53_7)*signed(FMAP_57_53);
			MULT_54(56)<=signed(DIN_54_7)*signed(FMAP_57_54);
			MULT_55(56)<=signed(DIN_55_7)*signed(FMAP_57_55);
			MULT_56(56)<=signed(DIN_56_7)*signed(FMAP_57_56);
			MULT_57(56)<=signed(DIN_57_7)*signed(FMAP_57_57);
			MULT_58(56)<=signed(DIN_58_7)*signed(FMAP_57_58);
			MULT_59(56)<=signed(DIN_59_7)*signed(FMAP_57_59);
			MULT_60(56)<=signed(DIN_60_7)*signed(FMAP_57_60);
			MULT_61(56)<=signed(DIN_61_7)*signed(FMAP_57_61);
			MULT_62(56)<=signed(DIN_62_7)*signed(FMAP_57_62);
			MULT_63(56)<=signed(DIN_63_7)*signed(FMAP_57_63);
			MULT_64(56)<=signed(DIN_64_7)*signed(FMAP_57_64);
			MULT_65(56)<=signed(DIN_65_7)*signed(FMAP_57_65);
			MULT_66(56)<=signed(DIN_66_7)*signed(FMAP_57_66);
			MULT_67(56)<=signed(DIN_67_7)*signed(FMAP_57_67);
			MULT_68(56)<=signed(DIN_68_7)*signed(FMAP_57_68);
			MULT_69(56)<=signed(DIN_69_7)*signed(FMAP_57_69);
			MULT_70(56)<=signed(DIN_70_7)*signed(FMAP_57_70);
			MULT_71(56)<=signed(DIN_71_7)*signed(FMAP_57_71);
			MULT_72(56)<=signed(DIN_72_7)*signed(FMAP_57_72);
			MULT_73(56)<=signed(DIN_73_7)*signed(FMAP_57_73);
			MULT_74(56)<=signed(DIN_74_7)*signed(FMAP_57_74);
			MULT_75(56)<=signed(DIN_75_7)*signed(FMAP_57_75);
			MULT_76(56)<=signed(DIN_76_7)*signed(FMAP_57_76);
			MULT_77(56)<=signed(DIN_77_7)*signed(FMAP_57_77);
			MULT_78(56)<=signed(DIN_78_7)*signed(FMAP_57_78);
			MULT_79(56)<=signed(DIN_79_7)*signed(FMAP_57_79);
			MULT_80(56)<=signed(DIN_80_7)*signed(FMAP_57_80);
			MULT_81(56)<=signed(DIN_81_7)*signed(FMAP_57_81);
			MULT_82(56)<=signed(DIN_82_7)*signed(FMAP_57_82);
			MULT_83(56)<=signed(DIN_83_7)*signed(FMAP_57_83);
			MULT_84(56)<=signed(DIN_84_7)*signed(FMAP_57_84);
			MULT_85(56)<=signed(DIN_85_7)*signed(FMAP_57_85);
			MULT_86(56)<=signed(DIN_86_7)*signed(FMAP_57_86);
			MULT_87(56)<=signed(DIN_87_7)*signed(FMAP_57_87);
			MULT_88(56)<=signed(DIN_88_7)*signed(FMAP_57_88);
			MULT_89(56)<=signed(DIN_89_7)*signed(FMAP_57_89);
			MULT_90(56)<=signed(DIN_90_7)*signed(FMAP_57_90);
			MULT_91(56)<=signed(DIN_91_7)*signed(FMAP_57_91);
			MULT_92(56)<=signed(DIN_92_7)*signed(FMAP_57_92);
			MULT_93(56)<=signed(DIN_93_7)*signed(FMAP_57_93);
			MULT_94(56)<=signed(DIN_94_7)*signed(FMAP_57_94);
			MULT_95(56)<=signed(DIN_95_7)*signed(FMAP_57_95);
			MULT_96(56)<=signed(DIN_96_7)*signed(FMAP_57_96);
			MULT_97(56)<=signed(DIN_97_7)*signed(FMAP_57_97);
			MULT_98(56)<=signed(DIN_98_7)*signed(FMAP_57_98);
			MULT_99(56)<=signed(DIN_99_7)*signed(FMAP_57_99);
			MULT_100(56)<=signed(DIN_100_7)*signed(FMAP_57_100);
			MULT_101(56)<=signed(DIN_101_7)*signed(FMAP_57_101);
			MULT_102(56)<=signed(DIN_102_7)*signed(FMAP_57_102);
			MULT_103(56)<=signed(DIN_103_7)*signed(FMAP_57_103);
			MULT_104(56)<=signed(DIN_104_7)*signed(FMAP_57_104);
			MULT_105(56)<=signed(DIN_105_7)*signed(FMAP_57_105);
			MULT_106(56)<=signed(DIN_106_7)*signed(FMAP_57_106);
			MULT_107(56)<=signed(DIN_107_7)*signed(FMAP_57_107);
			MULT_108(56)<=signed(DIN_108_7)*signed(FMAP_57_108);
			MULT_109(56)<=signed(DIN_109_7)*signed(FMAP_57_109);
			MULT_110(56)<=signed(DIN_110_7)*signed(FMAP_57_110);
			MULT_111(56)<=signed(DIN_111_7)*signed(FMAP_57_111);
			MULT_112(56)<=signed(DIN_112_7)*signed(FMAP_57_112);
			MULT_113(56)<=signed(DIN_113_7)*signed(FMAP_57_113);
			MULT_114(56)<=signed(DIN_114_7)*signed(FMAP_57_114);
			MULT_115(56)<=signed(DIN_115_7)*signed(FMAP_57_115);
			MULT_116(56)<=signed(DIN_116_7)*signed(FMAP_57_116);
			MULT_117(56)<=signed(DIN_117_7)*signed(FMAP_57_117);
			MULT_118(56)<=signed(DIN_118_7)*signed(FMAP_57_118);
			MULT_119(56)<=signed(DIN_119_7)*signed(FMAP_57_119);
			MULT_120(56)<=signed(DIN_120_7)*signed(FMAP_57_120);

			MULT_1(57)<=signed(DIN_1_7)*signed(FMAP_58_1);
			MULT_2(57)<=signed(DIN_2_7)*signed(FMAP_58_2);
			MULT_3(57)<=signed(DIN_3_7)*signed(FMAP_58_3);
			MULT_4(57)<=signed(DIN_4_7)*signed(FMAP_58_4);
			MULT_5(57)<=signed(DIN_5_7)*signed(FMAP_58_5);
			MULT_6(57)<=signed(DIN_6_7)*signed(FMAP_58_6);
			MULT_7(57)<=signed(DIN_7_7)*signed(FMAP_58_7);
			MULT_8(57)<=signed(DIN_8_7)*signed(FMAP_58_8);
			MULT_9(57)<=signed(DIN_9_7)*signed(FMAP_58_9);
			MULT_10(57)<=signed(DIN_10_7)*signed(FMAP_58_10);
			MULT_11(57)<=signed(DIN_11_7)*signed(FMAP_58_11);
			MULT_12(57)<=signed(DIN_12_7)*signed(FMAP_58_12);
			MULT_13(57)<=signed(DIN_13_7)*signed(FMAP_58_13);
			MULT_14(57)<=signed(DIN_14_7)*signed(FMAP_58_14);
			MULT_15(57)<=signed(DIN_15_7)*signed(FMAP_58_15);
			MULT_16(57)<=signed(DIN_16_7)*signed(FMAP_58_16);
			MULT_17(57)<=signed(DIN_17_7)*signed(FMAP_58_17);
			MULT_18(57)<=signed(DIN_18_7)*signed(FMAP_58_18);
			MULT_19(57)<=signed(DIN_19_7)*signed(FMAP_58_19);
			MULT_20(57)<=signed(DIN_20_7)*signed(FMAP_58_20);
			MULT_21(57)<=signed(DIN_21_7)*signed(FMAP_58_21);
			MULT_22(57)<=signed(DIN_22_7)*signed(FMAP_58_22);
			MULT_23(57)<=signed(DIN_23_7)*signed(FMAP_58_23);
			MULT_24(57)<=signed(DIN_24_7)*signed(FMAP_58_24);
			MULT_25(57)<=signed(DIN_25_7)*signed(FMAP_58_25);
			MULT_26(57)<=signed(DIN_26_7)*signed(FMAP_58_26);
			MULT_27(57)<=signed(DIN_27_7)*signed(FMAP_58_27);
			MULT_28(57)<=signed(DIN_28_7)*signed(FMAP_58_28);
			MULT_29(57)<=signed(DIN_29_7)*signed(FMAP_58_29);
			MULT_30(57)<=signed(DIN_30_7)*signed(FMAP_58_30);
			MULT_31(57)<=signed(DIN_31_7)*signed(FMAP_58_31);
			MULT_32(57)<=signed(DIN_32_7)*signed(FMAP_58_32);
			MULT_33(57)<=signed(DIN_33_7)*signed(FMAP_58_33);
			MULT_34(57)<=signed(DIN_34_7)*signed(FMAP_58_34);
			MULT_35(57)<=signed(DIN_35_7)*signed(FMAP_58_35);
			MULT_36(57)<=signed(DIN_36_7)*signed(FMAP_58_36);
			MULT_37(57)<=signed(DIN_37_7)*signed(FMAP_58_37);
			MULT_38(57)<=signed(DIN_38_7)*signed(FMAP_58_38);
			MULT_39(57)<=signed(DIN_39_7)*signed(FMAP_58_39);
			MULT_40(57)<=signed(DIN_40_7)*signed(FMAP_58_40);
			MULT_41(57)<=signed(DIN_41_7)*signed(FMAP_58_41);
			MULT_42(57)<=signed(DIN_42_7)*signed(FMAP_58_42);
			MULT_43(57)<=signed(DIN_43_7)*signed(FMAP_58_43);
			MULT_44(57)<=signed(DIN_44_7)*signed(FMAP_58_44);
			MULT_45(57)<=signed(DIN_45_7)*signed(FMAP_58_45);
			MULT_46(57)<=signed(DIN_46_7)*signed(FMAP_58_46);
			MULT_47(57)<=signed(DIN_47_7)*signed(FMAP_58_47);
			MULT_48(57)<=signed(DIN_48_7)*signed(FMAP_58_48);
			MULT_49(57)<=signed(DIN_49_7)*signed(FMAP_58_49);
			MULT_50(57)<=signed(DIN_50_7)*signed(FMAP_58_50);
			MULT_51(57)<=signed(DIN_51_7)*signed(FMAP_58_51);
			MULT_52(57)<=signed(DIN_52_7)*signed(FMAP_58_52);
			MULT_53(57)<=signed(DIN_53_7)*signed(FMAP_58_53);
			MULT_54(57)<=signed(DIN_54_7)*signed(FMAP_58_54);
			MULT_55(57)<=signed(DIN_55_7)*signed(FMAP_58_55);
			MULT_56(57)<=signed(DIN_56_7)*signed(FMAP_58_56);
			MULT_57(57)<=signed(DIN_57_7)*signed(FMAP_58_57);
			MULT_58(57)<=signed(DIN_58_7)*signed(FMAP_58_58);
			MULT_59(57)<=signed(DIN_59_7)*signed(FMAP_58_59);
			MULT_60(57)<=signed(DIN_60_7)*signed(FMAP_58_60);
			MULT_61(57)<=signed(DIN_61_7)*signed(FMAP_58_61);
			MULT_62(57)<=signed(DIN_62_7)*signed(FMAP_58_62);
			MULT_63(57)<=signed(DIN_63_7)*signed(FMAP_58_63);
			MULT_64(57)<=signed(DIN_64_7)*signed(FMAP_58_64);
			MULT_65(57)<=signed(DIN_65_7)*signed(FMAP_58_65);
			MULT_66(57)<=signed(DIN_66_7)*signed(FMAP_58_66);
			MULT_67(57)<=signed(DIN_67_7)*signed(FMAP_58_67);
			MULT_68(57)<=signed(DIN_68_7)*signed(FMAP_58_68);
			MULT_69(57)<=signed(DIN_69_7)*signed(FMAP_58_69);
			MULT_70(57)<=signed(DIN_70_7)*signed(FMAP_58_70);
			MULT_71(57)<=signed(DIN_71_7)*signed(FMAP_58_71);
			MULT_72(57)<=signed(DIN_72_7)*signed(FMAP_58_72);
			MULT_73(57)<=signed(DIN_73_7)*signed(FMAP_58_73);
			MULT_74(57)<=signed(DIN_74_7)*signed(FMAP_58_74);
			MULT_75(57)<=signed(DIN_75_7)*signed(FMAP_58_75);
			MULT_76(57)<=signed(DIN_76_7)*signed(FMAP_58_76);
			MULT_77(57)<=signed(DIN_77_7)*signed(FMAP_58_77);
			MULT_78(57)<=signed(DIN_78_7)*signed(FMAP_58_78);
			MULT_79(57)<=signed(DIN_79_7)*signed(FMAP_58_79);
			MULT_80(57)<=signed(DIN_80_7)*signed(FMAP_58_80);
			MULT_81(57)<=signed(DIN_81_7)*signed(FMAP_58_81);
			MULT_82(57)<=signed(DIN_82_7)*signed(FMAP_58_82);
			MULT_83(57)<=signed(DIN_83_7)*signed(FMAP_58_83);
			MULT_84(57)<=signed(DIN_84_7)*signed(FMAP_58_84);
			MULT_85(57)<=signed(DIN_85_7)*signed(FMAP_58_85);
			MULT_86(57)<=signed(DIN_86_7)*signed(FMAP_58_86);
			MULT_87(57)<=signed(DIN_87_7)*signed(FMAP_58_87);
			MULT_88(57)<=signed(DIN_88_7)*signed(FMAP_58_88);
			MULT_89(57)<=signed(DIN_89_7)*signed(FMAP_58_89);
			MULT_90(57)<=signed(DIN_90_7)*signed(FMAP_58_90);
			MULT_91(57)<=signed(DIN_91_7)*signed(FMAP_58_91);
			MULT_92(57)<=signed(DIN_92_7)*signed(FMAP_58_92);
			MULT_93(57)<=signed(DIN_93_7)*signed(FMAP_58_93);
			MULT_94(57)<=signed(DIN_94_7)*signed(FMAP_58_94);
			MULT_95(57)<=signed(DIN_95_7)*signed(FMAP_58_95);
			MULT_96(57)<=signed(DIN_96_7)*signed(FMAP_58_96);
			MULT_97(57)<=signed(DIN_97_7)*signed(FMAP_58_97);
			MULT_98(57)<=signed(DIN_98_7)*signed(FMAP_58_98);
			MULT_99(57)<=signed(DIN_99_7)*signed(FMAP_58_99);
			MULT_100(57)<=signed(DIN_100_7)*signed(FMAP_58_100);
			MULT_101(57)<=signed(DIN_101_7)*signed(FMAP_58_101);
			MULT_102(57)<=signed(DIN_102_7)*signed(FMAP_58_102);
			MULT_103(57)<=signed(DIN_103_7)*signed(FMAP_58_103);
			MULT_104(57)<=signed(DIN_104_7)*signed(FMAP_58_104);
			MULT_105(57)<=signed(DIN_105_7)*signed(FMAP_58_105);
			MULT_106(57)<=signed(DIN_106_7)*signed(FMAP_58_106);
			MULT_107(57)<=signed(DIN_107_7)*signed(FMAP_58_107);
			MULT_108(57)<=signed(DIN_108_7)*signed(FMAP_58_108);
			MULT_109(57)<=signed(DIN_109_7)*signed(FMAP_58_109);
			MULT_110(57)<=signed(DIN_110_7)*signed(FMAP_58_110);
			MULT_111(57)<=signed(DIN_111_7)*signed(FMAP_58_111);
			MULT_112(57)<=signed(DIN_112_7)*signed(FMAP_58_112);
			MULT_113(57)<=signed(DIN_113_7)*signed(FMAP_58_113);
			MULT_114(57)<=signed(DIN_114_7)*signed(FMAP_58_114);
			MULT_115(57)<=signed(DIN_115_7)*signed(FMAP_58_115);
			MULT_116(57)<=signed(DIN_116_7)*signed(FMAP_58_116);
			MULT_117(57)<=signed(DIN_117_7)*signed(FMAP_58_117);
			MULT_118(57)<=signed(DIN_118_7)*signed(FMAP_58_118);
			MULT_119(57)<=signed(DIN_119_7)*signed(FMAP_58_119);
			MULT_120(57)<=signed(DIN_120_7)*signed(FMAP_58_120);

			MULT_1(58)<=signed(DIN_1_7)*signed(FMAP_59_1);
			MULT_2(58)<=signed(DIN_2_7)*signed(FMAP_59_2);
			MULT_3(58)<=signed(DIN_3_7)*signed(FMAP_59_3);
			MULT_4(58)<=signed(DIN_4_7)*signed(FMAP_59_4);
			MULT_5(58)<=signed(DIN_5_7)*signed(FMAP_59_5);
			MULT_6(58)<=signed(DIN_6_7)*signed(FMAP_59_6);
			MULT_7(58)<=signed(DIN_7_7)*signed(FMAP_59_7);
			MULT_8(58)<=signed(DIN_8_7)*signed(FMAP_59_8);
			MULT_9(58)<=signed(DIN_9_7)*signed(FMAP_59_9);
			MULT_10(58)<=signed(DIN_10_7)*signed(FMAP_59_10);
			MULT_11(58)<=signed(DIN_11_7)*signed(FMAP_59_11);
			MULT_12(58)<=signed(DIN_12_7)*signed(FMAP_59_12);
			MULT_13(58)<=signed(DIN_13_7)*signed(FMAP_59_13);
			MULT_14(58)<=signed(DIN_14_7)*signed(FMAP_59_14);
			MULT_15(58)<=signed(DIN_15_7)*signed(FMAP_59_15);
			MULT_16(58)<=signed(DIN_16_7)*signed(FMAP_59_16);
			MULT_17(58)<=signed(DIN_17_7)*signed(FMAP_59_17);
			MULT_18(58)<=signed(DIN_18_7)*signed(FMAP_59_18);
			MULT_19(58)<=signed(DIN_19_7)*signed(FMAP_59_19);
			MULT_20(58)<=signed(DIN_20_7)*signed(FMAP_59_20);
			MULT_21(58)<=signed(DIN_21_7)*signed(FMAP_59_21);
			MULT_22(58)<=signed(DIN_22_7)*signed(FMAP_59_22);
			MULT_23(58)<=signed(DIN_23_7)*signed(FMAP_59_23);
			MULT_24(58)<=signed(DIN_24_7)*signed(FMAP_59_24);
			MULT_25(58)<=signed(DIN_25_7)*signed(FMAP_59_25);
			MULT_26(58)<=signed(DIN_26_7)*signed(FMAP_59_26);
			MULT_27(58)<=signed(DIN_27_7)*signed(FMAP_59_27);
			MULT_28(58)<=signed(DIN_28_7)*signed(FMAP_59_28);
			MULT_29(58)<=signed(DIN_29_7)*signed(FMAP_59_29);
			MULT_30(58)<=signed(DIN_30_7)*signed(FMAP_59_30);
			MULT_31(58)<=signed(DIN_31_7)*signed(FMAP_59_31);
			MULT_32(58)<=signed(DIN_32_7)*signed(FMAP_59_32);
			MULT_33(58)<=signed(DIN_33_7)*signed(FMAP_59_33);
			MULT_34(58)<=signed(DIN_34_7)*signed(FMAP_59_34);
			MULT_35(58)<=signed(DIN_35_7)*signed(FMAP_59_35);
			MULT_36(58)<=signed(DIN_36_7)*signed(FMAP_59_36);
			MULT_37(58)<=signed(DIN_37_7)*signed(FMAP_59_37);
			MULT_38(58)<=signed(DIN_38_7)*signed(FMAP_59_38);
			MULT_39(58)<=signed(DIN_39_7)*signed(FMAP_59_39);
			MULT_40(58)<=signed(DIN_40_7)*signed(FMAP_59_40);
			MULT_41(58)<=signed(DIN_41_7)*signed(FMAP_59_41);
			MULT_42(58)<=signed(DIN_42_7)*signed(FMAP_59_42);
			MULT_43(58)<=signed(DIN_43_7)*signed(FMAP_59_43);
			MULT_44(58)<=signed(DIN_44_7)*signed(FMAP_59_44);
			MULT_45(58)<=signed(DIN_45_7)*signed(FMAP_59_45);
			MULT_46(58)<=signed(DIN_46_7)*signed(FMAP_59_46);
			MULT_47(58)<=signed(DIN_47_7)*signed(FMAP_59_47);
			MULT_48(58)<=signed(DIN_48_7)*signed(FMAP_59_48);
			MULT_49(58)<=signed(DIN_49_7)*signed(FMAP_59_49);
			MULT_50(58)<=signed(DIN_50_7)*signed(FMAP_59_50);
			MULT_51(58)<=signed(DIN_51_7)*signed(FMAP_59_51);
			MULT_52(58)<=signed(DIN_52_7)*signed(FMAP_59_52);
			MULT_53(58)<=signed(DIN_53_7)*signed(FMAP_59_53);
			MULT_54(58)<=signed(DIN_54_7)*signed(FMAP_59_54);
			MULT_55(58)<=signed(DIN_55_7)*signed(FMAP_59_55);
			MULT_56(58)<=signed(DIN_56_7)*signed(FMAP_59_56);
			MULT_57(58)<=signed(DIN_57_7)*signed(FMAP_59_57);
			MULT_58(58)<=signed(DIN_58_7)*signed(FMAP_59_58);
			MULT_59(58)<=signed(DIN_59_7)*signed(FMAP_59_59);
			MULT_60(58)<=signed(DIN_60_7)*signed(FMAP_59_60);
			MULT_61(58)<=signed(DIN_61_7)*signed(FMAP_59_61);
			MULT_62(58)<=signed(DIN_62_7)*signed(FMAP_59_62);
			MULT_63(58)<=signed(DIN_63_7)*signed(FMAP_59_63);
			MULT_64(58)<=signed(DIN_64_7)*signed(FMAP_59_64);
			MULT_65(58)<=signed(DIN_65_7)*signed(FMAP_59_65);
			MULT_66(58)<=signed(DIN_66_7)*signed(FMAP_59_66);
			MULT_67(58)<=signed(DIN_67_7)*signed(FMAP_59_67);
			MULT_68(58)<=signed(DIN_68_7)*signed(FMAP_59_68);
			MULT_69(58)<=signed(DIN_69_7)*signed(FMAP_59_69);
			MULT_70(58)<=signed(DIN_70_7)*signed(FMAP_59_70);
			MULT_71(58)<=signed(DIN_71_7)*signed(FMAP_59_71);
			MULT_72(58)<=signed(DIN_72_7)*signed(FMAP_59_72);
			MULT_73(58)<=signed(DIN_73_7)*signed(FMAP_59_73);
			MULT_74(58)<=signed(DIN_74_7)*signed(FMAP_59_74);
			MULT_75(58)<=signed(DIN_75_7)*signed(FMAP_59_75);
			MULT_76(58)<=signed(DIN_76_7)*signed(FMAP_59_76);
			MULT_77(58)<=signed(DIN_77_7)*signed(FMAP_59_77);
			MULT_78(58)<=signed(DIN_78_7)*signed(FMAP_59_78);
			MULT_79(58)<=signed(DIN_79_7)*signed(FMAP_59_79);
			MULT_80(58)<=signed(DIN_80_7)*signed(FMAP_59_80);
			MULT_81(58)<=signed(DIN_81_7)*signed(FMAP_59_81);
			MULT_82(58)<=signed(DIN_82_7)*signed(FMAP_59_82);
			MULT_83(58)<=signed(DIN_83_7)*signed(FMAP_59_83);
			MULT_84(58)<=signed(DIN_84_7)*signed(FMAP_59_84);
			MULT_85(58)<=signed(DIN_85_7)*signed(FMAP_59_85);
			MULT_86(58)<=signed(DIN_86_7)*signed(FMAP_59_86);
			MULT_87(58)<=signed(DIN_87_7)*signed(FMAP_59_87);
			MULT_88(58)<=signed(DIN_88_7)*signed(FMAP_59_88);
			MULT_89(58)<=signed(DIN_89_7)*signed(FMAP_59_89);
			MULT_90(58)<=signed(DIN_90_7)*signed(FMAP_59_90);
			MULT_91(58)<=signed(DIN_91_7)*signed(FMAP_59_91);
			MULT_92(58)<=signed(DIN_92_7)*signed(FMAP_59_92);
			MULT_93(58)<=signed(DIN_93_7)*signed(FMAP_59_93);
			MULT_94(58)<=signed(DIN_94_7)*signed(FMAP_59_94);
			MULT_95(58)<=signed(DIN_95_7)*signed(FMAP_59_95);
			MULT_96(58)<=signed(DIN_96_7)*signed(FMAP_59_96);
			MULT_97(58)<=signed(DIN_97_7)*signed(FMAP_59_97);
			MULT_98(58)<=signed(DIN_98_7)*signed(FMAP_59_98);
			MULT_99(58)<=signed(DIN_99_7)*signed(FMAP_59_99);
			MULT_100(58)<=signed(DIN_100_7)*signed(FMAP_59_100);
			MULT_101(58)<=signed(DIN_101_7)*signed(FMAP_59_101);
			MULT_102(58)<=signed(DIN_102_7)*signed(FMAP_59_102);
			MULT_103(58)<=signed(DIN_103_7)*signed(FMAP_59_103);
			MULT_104(58)<=signed(DIN_104_7)*signed(FMAP_59_104);
			MULT_105(58)<=signed(DIN_105_7)*signed(FMAP_59_105);
			MULT_106(58)<=signed(DIN_106_7)*signed(FMAP_59_106);
			MULT_107(58)<=signed(DIN_107_7)*signed(FMAP_59_107);
			MULT_108(58)<=signed(DIN_108_7)*signed(FMAP_59_108);
			MULT_109(58)<=signed(DIN_109_7)*signed(FMAP_59_109);
			MULT_110(58)<=signed(DIN_110_7)*signed(FMAP_59_110);
			MULT_111(58)<=signed(DIN_111_7)*signed(FMAP_59_111);
			MULT_112(58)<=signed(DIN_112_7)*signed(FMAP_59_112);
			MULT_113(58)<=signed(DIN_113_7)*signed(FMAP_59_113);
			MULT_114(58)<=signed(DIN_114_7)*signed(FMAP_59_114);
			MULT_115(58)<=signed(DIN_115_7)*signed(FMAP_59_115);
			MULT_116(58)<=signed(DIN_116_7)*signed(FMAP_59_116);
			MULT_117(58)<=signed(DIN_117_7)*signed(FMAP_59_117);
			MULT_118(58)<=signed(DIN_118_7)*signed(FMAP_59_118);
			MULT_119(58)<=signed(DIN_119_7)*signed(FMAP_59_119);
			MULT_120(58)<=signed(DIN_120_7)*signed(FMAP_59_120);

			MULT_1(59)<=signed(DIN_1_7)*signed(FMAP_60_1);
			MULT_2(59)<=signed(DIN_2_7)*signed(FMAP_60_2);
			MULT_3(59)<=signed(DIN_3_7)*signed(FMAP_60_3);
			MULT_4(59)<=signed(DIN_4_7)*signed(FMAP_60_4);
			MULT_5(59)<=signed(DIN_5_7)*signed(FMAP_60_5);
			MULT_6(59)<=signed(DIN_6_7)*signed(FMAP_60_6);
			MULT_7(59)<=signed(DIN_7_7)*signed(FMAP_60_7);
			MULT_8(59)<=signed(DIN_8_7)*signed(FMAP_60_8);
			MULT_9(59)<=signed(DIN_9_7)*signed(FMAP_60_9);
			MULT_10(59)<=signed(DIN_10_7)*signed(FMAP_60_10);
			MULT_11(59)<=signed(DIN_11_7)*signed(FMAP_60_11);
			MULT_12(59)<=signed(DIN_12_7)*signed(FMAP_60_12);
			MULT_13(59)<=signed(DIN_13_7)*signed(FMAP_60_13);
			MULT_14(59)<=signed(DIN_14_7)*signed(FMAP_60_14);
			MULT_15(59)<=signed(DIN_15_7)*signed(FMAP_60_15);
			MULT_16(59)<=signed(DIN_16_7)*signed(FMAP_60_16);
			MULT_17(59)<=signed(DIN_17_7)*signed(FMAP_60_17);
			MULT_18(59)<=signed(DIN_18_7)*signed(FMAP_60_18);
			MULT_19(59)<=signed(DIN_19_7)*signed(FMAP_60_19);
			MULT_20(59)<=signed(DIN_20_7)*signed(FMAP_60_20);
			MULT_21(59)<=signed(DIN_21_7)*signed(FMAP_60_21);
			MULT_22(59)<=signed(DIN_22_7)*signed(FMAP_60_22);
			MULT_23(59)<=signed(DIN_23_7)*signed(FMAP_60_23);
			MULT_24(59)<=signed(DIN_24_7)*signed(FMAP_60_24);
			MULT_25(59)<=signed(DIN_25_7)*signed(FMAP_60_25);
			MULT_26(59)<=signed(DIN_26_7)*signed(FMAP_60_26);
			MULT_27(59)<=signed(DIN_27_7)*signed(FMAP_60_27);
			MULT_28(59)<=signed(DIN_28_7)*signed(FMAP_60_28);
			MULT_29(59)<=signed(DIN_29_7)*signed(FMAP_60_29);
			MULT_30(59)<=signed(DIN_30_7)*signed(FMAP_60_30);
			MULT_31(59)<=signed(DIN_31_7)*signed(FMAP_60_31);
			MULT_32(59)<=signed(DIN_32_7)*signed(FMAP_60_32);
			MULT_33(59)<=signed(DIN_33_7)*signed(FMAP_60_33);
			MULT_34(59)<=signed(DIN_34_7)*signed(FMAP_60_34);
			MULT_35(59)<=signed(DIN_35_7)*signed(FMAP_60_35);
			MULT_36(59)<=signed(DIN_36_7)*signed(FMAP_60_36);
			MULT_37(59)<=signed(DIN_37_7)*signed(FMAP_60_37);
			MULT_38(59)<=signed(DIN_38_7)*signed(FMAP_60_38);
			MULT_39(59)<=signed(DIN_39_7)*signed(FMAP_60_39);
			MULT_40(59)<=signed(DIN_40_7)*signed(FMAP_60_40);
			MULT_41(59)<=signed(DIN_41_7)*signed(FMAP_60_41);
			MULT_42(59)<=signed(DIN_42_7)*signed(FMAP_60_42);
			MULT_43(59)<=signed(DIN_43_7)*signed(FMAP_60_43);
			MULT_44(59)<=signed(DIN_44_7)*signed(FMAP_60_44);
			MULT_45(59)<=signed(DIN_45_7)*signed(FMAP_60_45);
			MULT_46(59)<=signed(DIN_46_7)*signed(FMAP_60_46);
			MULT_47(59)<=signed(DIN_47_7)*signed(FMAP_60_47);
			MULT_48(59)<=signed(DIN_48_7)*signed(FMAP_60_48);
			MULT_49(59)<=signed(DIN_49_7)*signed(FMAP_60_49);
			MULT_50(59)<=signed(DIN_50_7)*signed(FMAP_60_50);
			MULT_51(59)<=signed(DIN_51_7)*signed(FMAP_60_51);
			MULT_52(59)<=signed(DIN_52_7)*signed(FMAP_60_52);
			MULT_53(59)<=signed(DIN_53_7)*signed(FMAP_60_53);
			MULT_54(59)<=signed(DIN_54_7)*signed(FMAP_60_54);
			MULT_55(59)<=signed(DIN_55_7)*signed(FMAP_60_55);
			MULT_56(59)<=signed(DIN_56_7)*signed(FMAP_60_56);
			MULT_57(59)<=signed(DIN_57_7)*signed(FMAP_60_57);
			MULT_58(59)<=signed(DIN_58_7)*signed(FMAP_60_58);
			MULT_59(59)<=signed(DIN_59_7)*signed(FMAP_60_59);
			MULT_60(59)<=signed(DIN_60_7)*signed(FMAP_60_60);
			MULT_61(59)<=signed(DIN_61_7)*signed(FMAP_60_61);
			MULT_62(59)<=signed(DIN_62_7)*signed(FMAP_60_62);
			MULT_63(59)<=signed(DIN_63_7)*signed(FMAP_60_63);
			MULT_64(59)<=signed(DIN_64_7)*signed(FMAP_60_64);
			MULT_65(59)<=signed(DIN_65_7)*signed(FMAP_60_65);
			MULT_66(59)<=signed(DIN_66_7)*signed(FMAP_60_66);
			MULT_67(59)<=signed(DIN_67_7)*signed(FMAP_60_67);
			MULT_68(59)<=signed(DIN_68_7)*signed(FMAP_60_68);
			MULT_69(59)<=signed(DIN_69_7)*signed(FMAP_60_69);
			MULT_70(59)<=signed(DIN_70_7)*signed(FMAP_60_70);
			MULT_71(59)<=signed(DIN_71_7)*signed(FMAP_60_71);
			MULT_72(59)<=signed(DIN_72_7)*signed(FMAP_60_72);
			MULT_73(59)<=signed(DIN_73_7)*signed(FMAP_60_73);
			MULT_74(59)<=signed(DIN_74_7)*signed(FMAP_60_74);
			MULT_75(59)<=signed(DIN_75_7)*signed(FMAP_60_75);
			MULT_76(59)<=signed(DIN_76_7)*signed(FMAP_60_76);
			MULT_77(59)<=signed(DIN_77_7)*signed(FMAP_60_77);
			MULT_78(59)<=signed(DIN_78_7)*signed(FMAP_60_78);
			MULT_79(59)<=signed(DIN_79_7)*signed(FMAP_60_79);
			MULT_80(59)<=signed(DIN_80_7)*signed(FMAP_60_80);
			MULT_81(59)<=signed(DIN_81_7)*signed(FMAP_60_81);
			MULT_82(59)<=signed(DIN_82_7)*signed(FMAP_60_82);
			MULT_83(59)<=signed(DIN_83_7)*signed(FMAP_60_83);
			MULT_84(59)<=signed(DIN_84_7)*signed(FMAP_60_84);
			MULT_85(59)<=signed(DIN_85_7)*signed(FMAP_60_85);
			MULT_86(59)<=signed(DIN_86_7)*signed(FMAP_60_86);
			MULT_87(59)<=signed(DIN_87_7)*signed(FMAP_60_87);
			MULT_88(59)<=signed(DIN_88_7)*signed(FMAP_60_88);
			MULT_89(59)<=signed(DIN_89_7)*signed(FMAP_60_89);
			MULT_90(59)<=signed(DIN_90_7)*signed(FMAP_60_90);
			MULT_91(59)<=signed(DIN_91_7)*signed(FMAP_60_91);
			MULT_92(59)<=signed(DIN_92_7)*signed(FMAP_60_92);
			MULT_93(59)<=signed(DIN_93_7)*signed(FMAP_60_93);
			MULT_94(59)<=signed(DIN_94_7)*signed(FMAP_60_94);
			MULT_95(59)<=signed(DIN_95_7)*signed(FMAP_60_95);
			MULT_96(59)<=signed(DIN_96_7)*signed(FMAP_60_96);
			MULT_97(59)<=signed(DIN_97_7)*signed(FMAP_60_97);
			MULT_98(59)<=signed(DIN_98_7)*signed(FMAP_60_98);
			MULT_99(59)<=signed(DIN_99_7)*signed(FMAP_60_99);
			MULT_100(59)<=signed(DIN_100_7)*signed(FMAP_60_100);
			MULT_101(59)<=signed(DIN_101_7)*signed(FMAP_60_101);
			MULT_102(59)<=signed(DIN_102_7)*signed(FMAP_60_102);
			MULT_103(59)<=signed(DIN_103_7)*signed(FMAP_60_103);
			MULT_104(59)<=signed(DIN_104_7)*signed(FMAP_60_104);
			MULT_105(59)<=signed(DIN_105_7)*signed(FMAP_60_105);
			MULT_106(59)<=signed(DIN_106_7)*signed(FMAP_60_106);
			MULT_107(59)<=signed(DIN_107_7)*signed(FMAP_60_107);
			MULT_108(59)<=signed(DIN_108_7)*signed(FMAP_60_108);
			MULT_109(59)<=signed(DIN_109_7)*signed(FMAP_60_109);
			MULT_110(59)<=signed(DIN_110_7)*signed(FMAP_60_110);
			MULT_111(59)<=signed(DIN_111_7)*signed(FMAP_60_111);
			MULT_112(59)<=signed(DIN_112_7)*signed(FMAP_60_112);
			MULT_113(59)<=signed(DIN_113_7)*signed(FMAP_60_113);
			MULT_114(59)<=signed(DIN_114_7)*signed(FMAP_60_114);
			MULT_115(59)<=signed(DIN_115_7)*signed(FMAP_60_115);
			MULT_116(59)<=signed(DIN_116_7)*signed(FMAP_60_116);
			MULT_117(59)<=signed(DIN_117_7)*signed(FMAP_60_117);
			MULT_118(59)<=signed(DIN_118_7)*signed(FMAP_60_118);
			MULT_119(59)<=signed(DIN_119_7)*signed(FMAP_60_119);
			MULT_120(59)<=signed(DIN_120_7)*signed(FMAP_60_120);

			MULT_1(60)<=signed(DIN_1_7)*signed(FMAP_61_1);
			MULT_2(60)<=signed(DIN_2_7)*signed(FMAP_61_2);
			MULT_3(60)<=signed(DIN_3_7)*signed(FMAP_61_3);
			MULT_4(60)<=signed(DIN_4_7)*signed(FMAP_61_4);
			MULT_5(60)<=signed(DIN_5_7)*signed(FMAP_61_5);
			MULT_6(60)<=signed(DIN_6_7)*signed(FMAP_61_6);
			MULT_7(60)<=signed(DIN_7_7)*signed(FMAP_61_7);
			MULT_8(60)<=signed(DIN_8_7)*signed(FMAP_61_8);
			MULT_9(60)<=signed(DIN_9_7)*signed(FMAP_61_9);
			MULT_10(60)<=signed(DIN_10_7)*signed(FMAP_61_10);
			MULT_11(60)<=signed(DIN_11_7)*signed(FMAP_61_11);
			MULT_12(60)<=signed(DIN_12_7)*signed(FMAP_61_12);
			MULT_13(60)<=signed(DIN_13_7)*signed(FMAP_61_13);
			MULT_14(60)<=signed(DIN_14_7)*signed(FMAP_61_14);
			MULT_15(60)<=signed(DIN_15_7)*signed(FMAP_61_15);
			MULT_16(60)<=signed(DIN_16_7)*signed(FMAP_61_16);
			MULT_17(60)<=signed(DIN_17_7)*signed(FMAP_61_17);
			MULT_18(60)<=signed(DIN_18_7)*signed(FMAP_61_18);
			MULT_19(60)<=signed(DIN_19_7)*signed(FMAP_61_19);
			MULT_20(60)<=signed(DIN_20_7)*signed(FMAP_61_20);
			MULT_21(60)<=signed(DIN_21_7)*signed(FMAP_61_21);
			MULT_22(60)<=signed(DIN_22_7)*signed(FMAP_61_22);
			MULT_23(60)<=signed(DIN_23_7)*signed(FMAP_61_23);
			MULT_24(60)<=signed(DIN_24_7)*signed(FMAP_61_24);
			MULT_25(60)<=signed(DIN_25_7)*signed(FMAP_61_25);
			MULT_26(60)<=signed(DIN_26_7)*signed(FMAP_61_26);
			MULT_27(60)<=signed(DIN_27_7)*signed(FMAP_61_27);
			MULT_28(60)<=signed(DIN_28_7)*signed(FMAP_61_28);
			MULT_29(60)<=signed(DIN_29_7)*signed(FMAP_61_29);
			MULT_30(60)<=signed(DIN_30_7)*signed(FMAP_61_30);
			MULT_31(60)<=signed(DIN_31_7)*signed(FMAP_61_31);
			MULT_32(60)<=signed(DIN_32_7)*signed(FMAP_61_32);
			MULT_33(60)<=signed(DIN_33_7)*signed(FMAP_61_33);
			MULT_34(60)<=signed(DIN_34_7)*signed(FMAP_61_34);
			MULT_35(60)<=signed(DIN_35_7)*signed(FMAP_61_35);
			MULT_36(60)<=signed(DIN_36_7)*signed(FMAP_61_36);
			MULT_37(60)<=signed(DIN_37_7)*signed(FMAP_61_37);
			MULT_38(60)<=signed(DIN_38_7)*signed(FMAP_61_38);
			MULT_39(60)<=signed(DIN_39_7)*signed(FMAP_61_39);
			MULT_40(60)<=signed(DIN_40_7)*signed(FMAP_61_40);
			MULT_41(60)<=signed(DIN_41_7)*signed(FMAP_61_41);
			MULT_42(60)<=signed(DIN_42_7)*signed(FMAP_61_42);
			MULT_43(60)<=signed(DIN_43_7)*signed(FMAP_61_43);
			MULT_44(60)<=signed(DIN_44_7)*signed(FMAP_61_44);
			MULT_45(60)<=signed(DIN_45_7)*signed(FMAP_61_45);
			MULT_46(60)<=signed(DIN_46_7)*signed(FMAP_61_46);
			MULT_47(60)<=signed(DIN_47_7)*signed(FMAP_61_47);
			MULT_48(60)<=signed(DIN_48_7)*signed(FMAP_61_48);
			MULT_49(60)<=signed(DIN_49_7)*signed(FMAP_61_49);
			MULT_50(60)<=signed(DIN_50_7)*signed(FMAP_61_50);
			MULT_51(60)<=signed(DIN_51_7)*signed(FMAP_61_51);
			MULT_52(60)<=signed(DIN_52_7)*signed(FMAP_61_52);
			MULT_53(60)<=signed(DIN_53_7)*signed(FMAP_61_53);
			MULT_54(60)<=signed(DIN_54_7)*signed(FMAP_61_54);
			MULT_55(60)<=signed(DIN_55_7)*signed(FMAP_61_55);
			MULT_56(60)<=signed(DIN_56_7)*signed(FMAP_61_56);
			MULT_57(60)<=signed(DIN_57_7)*signed(FMAP_61_57);
			MULT_58(60)<=signed(DIN_58_7)*signed(FMAP_61_58);
			MULT_59(60)<=signed(DIN_59_7)*signed(FMAP_61_59);
			MULT_60(60)<=signed(DIN_60_7)*signed(FMAP_61_60);
			MULT_61(60)<=signed(DIN_61_7)*signed(FMAP_61_61);
			MULT_62(60)<=signed(DIN_62_7)*signed(FMAP_61_62);
			MULT_63(60)<=signed(DIN_63_7)*signed(FMAP_61_63);
			MULT_64(60)<=signed(DIN_64_7)*signed(FMAP_61_64);
			MULT_65(60)<=signed(DIN_65_7)*signed(FMAP_61_65);
			MULT_66(60)<=signed(DIN_66_7)*signed(FMAP_61_66);
			MULT_67(60)<=signed(DIN_67_7)*signed(FMAP_61_67);
			MULT_68(60)<=signed(DIN_68_7)*signed(FMAP_61_68);
			MULT_69(60)<=signed(DIN_69_7)*signed(FMAP_61_69);
			MULT_70(60)<=signed(DIN_70_7)*signed(FMAP_61_70);
			MULT_71(60)<=signed(DIN_71_7)*signed(FMAP_61_71);
			MULT_72(60)<=signed(DIN_72_7)*signed(FMAP_61_72);
			MULT_73(60)<=signed(DIN_73_7)*signed(FMAP_61_73);
			MULT_74(60)<=signed(DIN_74_7)*signed(FMAP_61_74);
			MULT_75(60)<=signed(DIN_75_7)*signed(FMAP_61_75);
			MULT_76(60)<=signed(DIN_76_7)*signed(FMAP_61_76);
			MULT_77(60)<=signed(DIN_77_7)*signed(FMAP_61_77);
			MULT_78(60)<=signed(DIN_78_7)*signed(FMAP_61_78);
			MULT_79(60)<=signed(DIN_79_7)*signed(FMAP_61_79);
			MULT_80(60)<=signed(DIN_80_7)*signed(FMAP_61_80);
			MULT_81(60)<=signed(DIN_81_7)*signed(FMAP_61_81);
			MULT_82(60)<=signed(DIN_82_7)*signed(FMAP_61_82);
			MULT_83(60)<=signed(DIN_83_7)*signed(FMAP_61_83);
			MULT_84(60)<=signed(DIN_84_7)*signed(FMAP_61_84);
			MULT_85(60)<=signed(DIN_85_7)*signed(FMAP_61_85);
			MULT_86(60)<=signed(DIN_86_7)*signed(FMAP_61_86);
			MULT_87(60)<=signed(DIN_87_7)*signed(FMAP_61_87);
			MULT_88(60)<=signed(DIN_88_7)*signed(FMAP_61_88);
			MULT_89(60)<=signed(DIN_89_7)*signed(FMAP_61_89);
			MULT_90(60)<=signed(DIN_90_7)*signed(FMAP_61_90);
			MULT_91(60)<=signed(DIN_91_7)*signed(FMAP_61_91);
			MULT_92(60)<=signed(DIN_92_7)*signed(FMAP_61_92);
			MULT_93(60)<=signed(DIN_93_7)*signed(FMAP_61_93);
			MULT_94(60)<=signed(DIN_94_7)*signed(FMAP_61_94);
			MULT_95(60)<=signed(DIN_95_7)*signed(FMAP_61_95);
			MULT_96(60)<=signed(DIN_96_7)*signed(FMAP_61_96);
			MULT_97(60)<=signed(DIN_97_7)*signed(FMAP_61_97);
			MULT_98(60)<=signed(DIN_98_7)*signed(FMAP_61_98);
			MULT_99(60)<=signed(DIN_99_7)*signed(FMAP_61_99);
			MULT_100(60)<=signed(DIN_100_7)*signed(FMAP_61_100);
			MULT_101(60)<=signed(DIN_101_7)*signed(FMAP_61_101);
			MULT_102(60)<=signed(DIN_102_7)*signed(FMAP_61_102);
			MULT_103(60)<=signed(DIN_103_7)*signed(FMAP_61_103);
			MULT_104(60)<=signed(DIN_104_7)*signed(FMAP_61_104);
			MULT_105(60)<=signed(DIN_105_7)*signed(FMAP_61_105);
			MULT_106(60)<=signed(DIN_106_7)*signed(FMAP_61_106);
			MULT_107(60)<=signed(DIN_107_7)*signed(FMAP_61_107);
			MULT_108(60)<=signed(DIN_108_7)*signed(FMAP_61_108);
			MULT_109(60)<=signed(DIN_109_7)*signed(FMAP_61_109);
			MULT_110(60)<=signed(DIN_110_7)*signed(FMAP_61_110);
			MULT_111(60)<=signed(DIN_111_7)*signed(FMAP_61_111);
			MULT_112(60)<=signed(DIN_112_7)*signed(FMAP_61_112);
			MULT_113(60)<=signed(DIN_113_7)*signed(FMAP_61_113);
			MULT_114(60)<=signed(DIN_114_7)*signed(FMAP_61_114);
			MULT_115(60)<=signed(DIN_115_7)*signed(FMAP_61_115);
			MULT_116(60)<=signed(DIN_116_7)*signed(FMAP_61_116);
			MULT_117(60)<=signed(DIN_117_7)*signed(FMAP_61_117);
			MULT_118(60)<=signed(DIN_118_7)*signed(FMAP_61_118);
			MULT_119(60)<=signed(DIN_119_7)*signed(FMAP_61_119);
			MULT_120(60)<=signed(DIN_120_7)*signed(FMAP_61_120);

			MULT_1(61)<=signed(DIN_1_7)*signed(FMAP_62_1);
			MULT_2(61)<=signed(DIN_2_7)*signed(FMAP_62_2);
			MULT_3(61)<=signed(DIN_3_7)*signed(FMAP_62_3);
			MULT_4(61)<=signed(DIN_4_7)*signed(FMAP_62_4);
			MULT_5(61)<=signed(DIN_5_7)*signed(FMAP_62_5);
			MULT_6(61)<=signed(DIN_6_7)*signed(FMAP_62_6);
			MULT_7(61)<=signed(DIN_7_7)*signed(FMAP_62_7);
			MULT_8(61)<=signed(DIN_8_7)*signed(FMAP_62_8);
			MULT_9(61)<=signed(DIN_9_7)*signed(FMAP_62_9);
			MULT_10(61)<=signed(DIN_10_7)*signed(FMAP_62_10);
			MULT_11(61)<=signed(DIN_11_7)*signed(FMAP_62_11);
			MULT_12(61)<=signed(DIN_12_7)*signed(FMAP_62_12);
			MULT_13(61)<=signed(DIN_13_7)*signed(FMAP_62_13);
			MULT_14(61)<=signed(DIN_14_7)*signed(FMAP_62_14);
			MULT_15(61)<=signed(DIN_15_7)*signed(FMAP_62_15);
			MULT_16(61)<=signed(DIN_16_7)*signed(FMAP_62_16);
			MULT_17(61)<=signed(DIN_17_7)*signed(FMAP_62_17);
			MULT_18(61)<=signed(DIN_18_7)*signed(FMAP_62_18);
			MULT_19(61)<=signed(DIN_19_7)*signed(FMAP_62_19);
			MULT_20(61)<=signed(DIN_20_7)*signed(FMAP_62_20);
			MULT_21(61)<=signed(DIN_21_7)*signed(FMAP_62_21);
			MULT_22(61)<=signed(DIN_22_7)*signed(FMAP_62_22);
			MULT_23(61)<=signed(DIN_23_7)*signed(FMAP_62_23);
			MULT_24(61)<=signed(DIN_24_7)*signed(FMAP_62_24);
			MULT_25(61)<=signed(DIN_25_7)*signed(FMAP_62_25);
			MULT_26(61)<=signed(DIN_26_7)*signed(FMAP_62_26);
			MULT_27(61)<=signed(DIN_27_7)*signed(FMAP_62_27);
			MULT_28(61)<=signed(DIN_28_7)*signed(FMAP_62_28);
			MULT_29(61)<=signed(DIN_29_7)*signed(FMAP_62_29);
			MULT_30(61)<=signed(DIN_30_7)*signed(FMAP_62_30);
			MULT_31(61)<=signed(DIN_31_7)*signed(FMAP_62_31);
			MULT_32(61)<=signed(DIN_32_7)*signed(FMAP_62_32);
			MULT_33(61)<=signed(DIN_33_7)*signed(FMAP_62_33);
			MULT_34(61)<=signed(DIN_34_7)*signed(FMAP_62_34);
			MULT_35(61)<=signed(DIN_35_7)*signed(FMAP_62_35);
			MULT_36(61)<=signed(DIN_36_7)*signed(FMAP_62_36);
			MULT_37(61)<=signed(DIN_37_7)*signed(FMAP_62_37);
			MULT_38(61)<=signed(DIN_38_7)*signed(FMAP_62_38);
			MULT_39(61)<=signed(DIN_39_7)*signed(FMAP_62_39);
			MULT_40(61)<=signed(DIN_40_7)*signed(FMAP_62_40);
			MULT_41(61)<=signed(DIN_41_7)*signed(FMAP_62_41);
			MULT_42(61)<=signed(DIN_42_7)*signed(FMAP_62_42);
			MULT_43(61)<=signed(DIN_43_7)*signed(FMAP_62_43);
			MULT_44(61)<=signed(DIN_44_7)*signed(FMAP_62_44);
			MULT_45(61)<=signed(DIN_45_7)*signed(FMAP_62_45);
			MULT_46(61)<=signed(DIN_46_7)*signed(FMAP_62_46);
			MULT_47(61)<=signed(DIN_47_7)*signed(FMAP_62_47);
			MULT_48(61)<=signed(DIN_48_7)*signed(FMAP_62_48);
			MULT_49(61)<=signed(DIN_49_7)*signed(FMAP_62_49);
			MULT_50(61)<=signed(DIN_50_7)*signed(FMAP_62_50);
			MULT_51(61)<=signed(DIN_51_7)*signed(FMAP_62_51);
			MULT_52(61)<=signed(DIN_52_7)*signed(FMAP_62_52);
			MULT_53(61)<=signed(DIN_53_7)*signed(FMAP_62_53);
			MULT_54(61)<=signed(DIN_54_7)*signed(FMAP_62_54);
			MULT_55(61)<=signed(DIN_55_7)*signed(FMAP_62_55);
			MULT_56(61)<=signed(DIN_56_7)*signed(FMAP_62_56);
			MULT_57(61)<=signed(DIN_57_7)*signed(FMAP_62_57);
			MULT_58(61)<=signed(DIN_58_7)*signed(FMAP_62_58);
			MULT_59(61)<=signed(DIN_59_7)*signed(FMAP_62_59);
			MULT_60(61)<=signed(DIN_60_7)*signed(FMAP_62_60);
			MULT_61(61)<=signed(DIN_61_7)*signed(FMAP_62_61);
			MULT_62(61)<=signed(DIN_62_7)*signed(FMAP_62_62);
			MULT_63(61)<=signed(DIN_63_7)*signed(FMAP_62_63);
			MULT_64(61)<=signed(DIN_64_7)*signed(FMAP_62_64);
			MULT_65(61)<=signed(DIN_65_7)*signed(FMAP_62_65);
			MULT_66(61)<=signed(DIN_66_7)*signed(FMAP_62_66);
			MULT_67(61)<=signed(DIN_67_7)*signed(FMAP_62_67);
			MULT_68(61)<=signed(DIN_68_7)*signed(FMAP_62_68);
			MULT_69(61)<=signed(DIN_69_7)*signed(FMAP_62_69);
			MULT_70(61)<=signed(DIN_70_7)*signed(FMAP_62_70);
			MULT_71(61)<=signed(DIN_71_7)*signed(FMAP_62_71);
			MULT_72(61)<=signed(DIN_72_7)*signed(FMAP_62_72);
			MULT_73(61)<=signed(DIN_73_7)*signed(FMAP_62_73);
			MULT_74(61)<=signed(DIN_74_7)*signed(FMAP_62_74);
			MULT_75(61)<=signed(DIN_75_7)*signed(FMAP_62_75);
			MULT_76(61)<=signed(DIN_76_7)*signed(FMAP_62_76);
			MULT_77(61)<=signed(DIN_77_7)*signed(FMAP_62_77);
			MULT_78(61)<=signed(DIN_78_7)*signed(FMAP_62_78);
			MULT_79(61)<=signed(DIN_79_7)*signed(FMAP_62_79);
			MULT_80(61)<=signed(DIN_80_7)*signed(FMAP_62_80);
			MULT_81(61)<=signed(DIN_81_7)*signed(FMAP_62_81);
			MULT_82(61)<=signed(DIN_82_7)*signed(FMAP_62_82);
			MULT_83(61)<=signed(DIN_83_7)*signed(FMAP_62_83);
			MULT_84(61)<=signed(DIN_84_7)*signed(FMAP_62_84);
			MULT_85(61)<=signed(DIN_85_7)*signed(FMAP_62_85);
			MULT_86(61)<=signed(DIN_86_7)*signed(FMAP_62_86);
			MULT_87(61)<=signed(DIN_87_7)*signed(FMAP_62_87);
			MULT_88(61)<=signed(DIN_88_7)*signed(FMAP_62_88);
			MULT_89(61)<=signed(DIN_89_7)*signed(FMAP_62_89);
			MULT_90(61)<=signed(DIN_90_7)*signed(FMAP_62_90);
			MULT_91(61)<=signed(DIN_91_7)*signed(FMAP_62_91);
			MULT_92(61)<=signed(DIN_92_7)*signed(FMAP_62_92);
			MULT_93(61)<=signed(DIN_93_7)*signed(FMAP_62_93);
			MULT_94(61)<=signed(DIN_94_7)*signed(FMAP_62_94);
			MULT_95(61)<=signed(DIN_95_7)*signed(FMAP_62_95);
			MULT_96(61)<=signed(DIN_96_7)*signed(FMAP_62_96);
			MULT_97(61)<=signed(DIN_97_7)*signed(FMAP_62_97);
			MULT_98(61)<=signed(DIN_98_7)*signed(FMAP_62_98);
			MULT_99(61)<=signed(DIN_99_7)*signed(FMAP_62_99);
			MULT_100(61)<=signed(DIN_100_7)*signed(FMAP_62_100);
			MULT_101(61)<=signed(DIN_101_7)*signed(FMAP_62_101);
			MULT_102(61)<=signed(DIN_102_7)*signed(FMAP_62_102);
			MULT_103(61)<=signed(DIN_103_7)*signed(FMAP_62_103);
			MULT_104(61)<=signed(DIN_104_7)*signed(FMAP_62_104);
			MULT_105(61)<=signed(DIN_105_7)*signed(FMAP_62_105);
			MULT_106(61)<=signed(DIN_106_7)*signed(FMAP_62_106);
			MULT_107(61)<=signed(DIN_107_7)*signed(FMAP_62_107);
			MULT_108(61)<=signed(DIN_108_7)*signed(FMAP_62_108);
			MULT_109(61)<=signed(DIN_109_7)*signed(FMAP_62_109);
			MULT_110(61)<=signed(DIN_110_7)*signed(FMAP_62_110);
			MULT_111(61)<=signed(DIN_111_7)*signed(FMAP_62_111);
			MULT_112(61)<=signed(DIN_112_7)*signed(FMAP_62_112);
			MULT_113(61)<=signed(DIN_113_7)*signed(FMAP_62_113);
			MULT_114(61)<=signed(DIN_114_7)*signed(FMAP_62_114);
			MULT_115(61)<=signed(DIN_115_7)*signed(FMAP_62_115);
			MULT_116(61)<=signed(DIN_116_7)*signed(FMAP_62_116);
			MULT_117(61)<=signed(DIN_117_7)*signed(FMAP_62_117);
			MULT_118(61)<=signed(DIN_118_7)*signed(FMAP_62_118);
			MULT_119(61)<=signed(DIN_119_7)*signed(FMAP_62_119);
			MULT_120(61)<=signed(DIN_120_7)*signed(FMAP_62_120);

			MULT_1(62)<=signed(DIN_1_7)*signed(FMAP_63_1);
			MULT_2(62)<=signed(DIN_2_7)*signed(FMAP_63_2);
			MULT_3(62)<=signed(DIN_3_7)*signed(FMAP_63_3);
			MULT_4(62)<=signed(DIN_4_7)*signed(FMAP_63_4);
			MULT_5(62)<=signed(DIN_5_7)*signed(FMAP_63_5);
			MULT_6(62)<=signed(DIN_6_7)*signed(FMAP_63_6);
			MULT_7(62)<=signed(DIN_7_7)*signed(FMAP_63_7);
			MULT_8(62)<=signed(DIN_8_7)*signed(FMAP_63_8);
			MULT_9(62)<=signed(DIN_9_7)*signed(FMAP_63_9);
			MULT_10(62)<=signed(DIN_10_7)*signed(FMAP_63_10);
			MULT_11(62)<=signed(DIN_11_7)*signed(FMAP_63_11);
			MULT_12(62)<=signed(DIN_12_7)*signed(FMAP_63_12);
			MULT_13(62)<=signed(DIN_13_7)*signed(FMAP_63_13);
			MULT_14(62)<=signed(DIN_14_7)*signed(FMAP_63_14);
			MULT_15(62)<=signed(DIN_15_7)*signed(FMAP_63_15);
			MULT_16(62)<=signed(DIN_16_7)*signed(FMAP_63_16);
			MULT_17(62)<=signed(DIN_17_7)*signed(FMAP_63_17);
			MULT_18(62)<=signed(DIN_18_7)*signed(FMAP_63_18);
			MULT_19(62)<=signed(DIN_19_7)*signed(FMAP_63_19);
			MULT_20(62)<=signed(DIN_20_7)*signed(FMAP_63_20);
			MULT_21(62)<=signed(DIN_21_7)*signed(FMAP_63_21);
			MULT_22(62)<=signed(DIN_22_7)*signed(FMAP_63_22);
			MULT_23(62)<=signed(DIN_23_7)*signed(FMAP_63_23);
			MULT_24(62)<=signed(DIN_24_7)*signed(FMAP_63_24);
			MULT_25(62)<=signed(DIN_25_7)*signed(FMAP_63_25);
			MULT_26(62)<=signed(DIN_26_7)*signed(FMAP_63_26);
			MULT_27(62)<=signed(DIN_27_7)*signed(FMAP_63_27);
			MULT_28(62)<=signed(DIN_28_7)*signed(FMAP_63_28);
			MULT_29(62)<=signed(DIN_29_7)*signed(FMAP_63_29);
			MULT_30(62)<=signed(DIN_30_7)*signed(FMAP_63_30);
			MULT_31(62)<=signed(DIN_31_7)*signed(FMAP_63_31);
			MULT_32(62)<=signed(DIN_32_7)*signed(FMAP_63_32);
			MULT_33(62)<=signed(DIN_33_7)*signed(FMAP_63_33);
			MULT_34(62)<=signed(DIN_34_7)*signed(FMAP_63_34);
			MULT_35(62)<=signed(DIN_35_7)*signed(FMAP_63_35);
			MULT_36(62)<=signed(DIN_36_7)*signed(FMAP_63_36);
			MULT_37(62)<=signed(DIN_37_7)*signed(FMAP_63_37);
			MULT_38(62)<=signed(DIN_38_7)*signed(FMAP_63_38);
			MULT_39(62)<=signed(DIN_39_7)*signed(FMAP_63_39);
			MULT_40(62)<=signed(DIN_40_7)*signed(FMAP_63_40);
			MULT_41(62)<=signed(DIN_41_7)*signed(FMAP_63_41);
			MULT_42(62)<=signed(DIN_42_7)*signed(FMAP_63_42);
			MULT_43(62)<=signed(DIN_43_7)*signed(FMAP_63_43);
			MULT_44(62)<=signed(DIN_44_7)*signed(FMAP_63_44);
			MULT_45(62)<=signed(DIN_45_7)*signed(FMAP_63_45);
			MULT_46(62)<=signed(DIN_46_7)*signed(FMAP_63_46);
			MULT_47(62)<=signed(DIN_47_7)*signed(FMAP_63_47);
			MULT_48(62)<=signed(DIN_48_7)*signed(FMAP_63_48);
			MULT_49(62)<=signed(DIN_49_7)*signed(FMAP_63_49);
			MULT_50(62)<=signed(DIN_50_7)*signed(FMAP_63_50);
			MULT_51(62)<=signed(DIN_51_7)*signed(FMAP_63_51);
			MULT_52(62)<=signed(DIN_52_7)*signed(FMAP_63_52);
			MULT_53(62)<=signed(DIN_53_7)*signed(FMAP_63_53);
			MULT_54(62)<=signed(DIN_54_7)*signed(FMAP_63_54);
			MULT_55(62)<=signed(DIN_55_7)*signed(FMAP_63_55);
			MULT_56(62)<=signed(DIN_56_7)*signed(FMAP_63_56);
			MULT_57(62)<=signed(DIN_57_7)*signed(FMAP_63_57);
			MULT_58(62)<=signed(DIN_58_7)*signed(FMAP_63_58);
			MULT_59(62)<=signed(DIN_59_7)*signed(FMAP_63_59);
			MULT_60(62)<=signed(DIN_60_7)*signed(FMAP_63_60);
			MULT_61(62)<=signed(DIN_61_7)*signed(FMAP_63_61);
			MULT_62(62)<=signed(DIN_62_7)*signed(FMAP_63_62);
			MULT_63(62)<=signed(DIN_63_7)*signed(FMAP_63_63);
			MULT_64(62)<=signed(DIN_64_7)*signed(FMAP_63_64);
			MULT_65(62)<=signed(DIN_65_7)*signed(FMAP_63_65);
			MULT_66(62)<=signed(DIN_66_7)*signed(FMAP_63_66);
			MULT_67(62)<=signed(DIN_67_7)*signed(FMAP_63_67);
			MULT_68(62)<=signed(DIN_68_7)*signed(FMAP_63_68);
			MULT_69(62)<=signed(DIN_69_7)*signed(FMAP_63_69);
			MULT_70(62)<=signed(DIN_70_7)*signed(FMAP_63_70);
			MULT_71(62)<=signed(DIN_71_7)*signed(FMAP_63_71);
			MULT_72(62)<=signed(DIN_72_7)*signed(FMAP_63_72);
			MULT_73(62)<=signed(DIN_73_7)*signed(FMAP_63_73);
			MULT_74(62)<=signed(DIN_74_7)*signed(FMAP_63_74);
			MULT_75(62)<=signed(DIN_75_7)*signed(FMAP_63_75);
			MULT_76(62)<=signed(DIN_76_7)*signed(FMAP_63_76);
			MULT_77(62)<=signed(DIN_77_7)*signed(FMAP_63_77);
			MULT_78(62)<=signed(DIN_78_7)*signed(FMAP_63_78);
			MULT_79(62)<=signed(DIN_79_7)*signed(FMAP_63_79);
			MULT_80(62)<=signed(DIN_80_7)*signed(FMAP_63_80);
			MULT_81(62)<=signed(DIN_81_7)*signed(FMAP_63_81);
			MULT_82(62)<=signed(DIN_82_7)*signed(FMAP_63_82);
			MULT_83(62)<=signed(DIN_83_7)*signed(FMAP_63_83);
			MULT_84(62)<=signed(DIN_84_7)*signed(FMAP_63_84);
			MULT_85(62)<=signed(DIN_85_7)*signed(FMAP_63_85);
			MULT_86(62)<=signed(DIN_86_7)*signed(FMAP_63_86);
			MULT_87(62)<=signed(DIN_87_7)*signed(FMAP_63_87);
			MULT_88(62)<=signed(DIN_88_7)*signed(FMAP_63_88);
			MULT_89(62)<=signed(DIN_89_7)*signed(FMAP_63_89);
			MULT_90(62)<=signed(DIN_90_7)*signed(FMAP_63_90);
			MULT_91(62)<=signed(DIN_91_7)*signed(FMAP_63_91);
			MULT_92(62)<=signed(DIN_92_7)*signed(FMAP_63_92);
			MULT_93(62)<=signed(DIN_93_7)*signed(FMAP_63_93);
			MULT_94(62)<=signed(DIN_94_7)*signed(FMAP_63_94);
			MULT_95(62)<=signed(DIN_95_7)*signed(FMAP_63_95);
			MULT_96(62)<=signed(DIN_96_7)*signed(FMAP_63_96);
			MULT_97(62)<=signed(DIN_97_7)*signed(FMAP_63_97);
			MULT_98(62)<=signed(DIN_98_7)*signed(FMAP_63_98);
			MULT_99(62)<=signed(DIN_99_7)*signed(FMAP_63_99);
			MULT_100(62)<=signed(DIN_100_7)*signed(FMAP_63_100);
			MULT_101(62)<=signed(DIN_101_7)*signed(FMAP_63_101);
			MULT_102(62)<=signed(DIN_102_7)*signed(FMAP_63_102);
			MULT_103(62)<=signed(DIN_103_7)*signed(FMAP_63_103);
			MULT_104(62)<=signed(DIN_104_7)*signed(FMAP_63_104);
			MULT_105(62)<=signed(DIN_105_7)*signed(FMAP_63_105);
			MULT_106(62)<=signed(DIN_106_7)*signed(FMAP_63_106);
			MULT_107(62)<=signed(DIN_107_7)*signed(FMAP_63_107);
			MULT_108(62)<=signed(DIN_108_7)*signed(FMAP_63_108);
			MULT_109(62)<=signed(DIN_109_7)*signed(FMAP_63_109);
			MULT_110(62)<=signed(DIN_110_7)*signed(FMAP_63_110);
			MULT_111(62)<=signed(DIN_111_7)*signed(FMAP_63_111);
			MULT_112(62)<=signed(DIN_112_7)*signed(FMAP_63_112);
			MULT_113(62)<=signed(DIN_113_7)*signed(FMAP_63_113);
			MULT_114(62)<=signed(DIN_114_7)*signed(FMAP_63_114);
			MULT_115(62)<=signed(DIN_115_7)*signed(FMAP_63_115);
			MULT_116(62)<=signed(DIN_116_7)*signed(FMAP_63_116);
			MULT_117(62)<=signed(DIN_117_7)*signed(FMAP_63_117);
			MULT_118(62)<=signed(DIN_118_7)*signed(FMAP_63_118);
			MULT_119(62)<=signed(DIN_119_7)*signed(FMAP_63_119);
			MULT_120(62)<=signed(DIN_120_7)*signed(FMAP_63_120);

			MULT_1(63)<=signed(DIN_1_7)*signed(FMAP_64_1);
			MULT_2(63)<=signed(DIN_2_7)*signed(FMAP_64_2);
			MULT_3(63)<=signed(DIN_3_7)*signed(FMAP_64_3);
			MULT_4(63)<=signed(DIN_4_7)*signed(FMAP_64_4);
			MULT_5(63)<=signed(DIN_5_7)*signed(FMAP_64_5);
			MULT_6(63)<=signed(DIN_6_7)*signed(FMAP_64_6);
			MULT_7(63)<=signed(DIN_7_7)*signed(FMAP_64_7);
			MULT_8(63)<=signed(DIN_8_7)*signed(FMAP_64_8);
			MULT_9(63)<=signed(DIN_9_7)*signed(FMAP_64_9);
			MULT_10(63)<=signed(DIN_10_7)*signed(FMAP_64_10);
			MULT_11(63)<=signed(DIN_11_7)*signed(FMAP_64_11);
			MULT_12(63)<=signed(DIN_12_7)*signed(FMAP_64_12);
			MULT_13(63)<=signed(DIN_13_7)*signed(FMAP_64_13);
			MULT_14(63)<=signed(DIN_14_7)*signed(FMAP_64_14);
			MULT_15(63)<=signed(DIN_15_7)*signed(FMAP_64_15);
			MULT_16(63)<=signed(DIN_16_7)*signed(FMAP_64_16);
			MULT_17(63)<=signed(DIN_17_7)*signed(FMAP_64_17);
			MULT_18(63)<=signed(DIN_18_7)*signed(FMAP_64_18);
			MULT_19(63)<=signed(DIN_19_7)*signed(FMAP_64_19);
			MULT_20(63)<=signed(DIN_20_7)*signed(FMAP_64_20);
			MULT_21(63)<=signed(DIN_21_7)*signed(FMAP_64_21);
			MULT_22(63)<=signed(DIN_22_7)*signed(FMAP_64_22);
			MULT_23(63)<=signed(DIN_23_7)*signed(FMAP_64_23);
			MULT_24(63)<=signed(DIN_24_7)*signed(FMAP_64_24);
			MULT_25(63)<=signed(DIN_25_7)*signed(FMAP_64_25);
			MULT_26(63)<=signed(DIN_26_7)*signed(FMAP_64_26);
			MULT_27(63)<=signed(DIN_27_7)*signed(FMAP_64_27);
			MULT_28(63)<=signed(DIN_28_7)*signed(FMAP_64_28);
			MULT_29(63)<=signed(DIN_29_7)*signed(FMAP_64_29);
			MULT_30(63)<=signed(DIN_30_7)*signed(FMAP_64_30);
			MULT_31(63)<=signed(DIN_31_7)*signed(FMAP_64_31);
			MULT_32(63)<=signed(DIN_32_7)*signed(FMAP_64_32);
			MULT_33(63)<=signed(DIN_33_7)*signed(FMAP_64_33);
			MULT_34(63)<=signed(DIN_34_7)*signed(FMAP_64_34);
			MULT_35(63)<=signed(DIN_35_7)*signed(FMAP_64_35);
			MULT_36(63)<=signed(DIN_36_7)*signed(FMAP_64_36);
			MULT_37(63)<=signed(DIN_37_7)*signed(FMAP_64_37);
			MULT_38(63)<=signed(DIN_38_7)*signed(FMAP_64_38);
			MULT_39(63)<=signed(DIN_39_7)*signed(FMAP_64_39);
			MULT_40(63)<=signed(DIN_40_7)*signed(FMAP_64_40);
			MULT_41(63)<=signed(DIN_41_7)*signed(FMAP_64_41);
			MULT_42(63)<=signed(DIN_42_7)*signed(FMAP_64_42);
			MULT_43(63)<=signed(DIN_43_7)*signed(FMAP_64_43);
			MULT_44(63)<=signed(DIN_44_7)*signed(FMAP_64_44);
			MULT_45(63)<=signed(DIN_45_7)*signed(FMAP_64_45);
			MULT_46(63)<=signed(DIN_46_7)*signed(FMAP_64_46);
			MULT_47(63)<=signed(DIN_47_7)*signed(FMAP_64_47);
			MULT_48(63)<=signed(DIN_48_7)*signed(FMAP_64_48);
			MULT_49(63)<=signed(DIN_49_7)*signed(FMAP_64_49);
			MULT_50(63)<=signed(DIN_50_7)*signed(FMAP_64_50);
			MULT_51(63)<=signed(DIN_51_7)*signed(FMAP_64_51);
			MULT_52(63)<=signed(DIN_52_7)*signed(FMAP_64_52);
			MULT_53(63)<=signed(DIN_53_7)*signed(FMAP_64_53);
			MULT_54(63)<=signed(DIN_54_7)*signed(FMAP_64_54);
			MULT_55(63)<=signed(DIN_55_7)*signed(FMAP_64_55);
			MULT_56(63)<=signed(DIN_56_7)*signed(FMAP_64_56);
			MULT_57(63)<=signed(DIN_57_7)*signed(FMAP_64_57);
			MULT_58(63)<=signed(DIN_58_7)*signed(FMAP_64_58);
			MULT_59(63)<=signed(DIN_59_7)*signed(FMAP_64_59);
			MULT_60(63)<=signed(DIN_60_7)*signed(FMAP_64_60);
			MULT_61(63)<=signed(DIN_61_7)*signed(FMAP_64_61);
			MULT_62(63)<=signed(DIN_62_7)*signed(FMAP_64_62);
			MULT_63(63)<=signed(DIN_63_7)*signed(FMAP_64_63);
			MULT_64(63)<=signed(DIN_64_7)*signed(FMAP_64_64);
			MULT_65(63)<=signed(DIN_65_7)*signed(FMAP_64_65);
			MULT_66(63)<=signed(DIN_66_7)*signed(FMAP_64_66);
			MULT_67(63)<=signed(DIN_67_7)*signed(FMAP_64_67);
			MULT_68(63)<=signed(DIN_68_7)*signed(FMAP_64_68);
			MULT_69(63)<=signed(DIN_69_7)*signed(FMAP_64_69);
			MULT_70(63)<=signed(DIN_70_7)*signed(FMAP_64_70);
			MULT_71(63)<=signed(DIN_71_7)*signed(FMAP_64_71);
			MULT_72(63)<=signed(DIN_72_7)*signed(FMAP_64_72);
			MULT_73(63)<=signed(DIN_73_7)*signed(FMAP_64_73);
			MULT_74(63)<=signed(DIN_74_7)*signed(FMAP_64_74);
			MULT_75(63)<=signed(DIN_75_7)*signed(FMAP_64_75);
			MULT_76(63)<=signed(DIN_76_7)*signed(FMAP_64_76);
			MULT_77(63)<=signed(DIN_77_7)*signed(FMAP_64_77);
			MULT_78(63)<=signed(DIN_78_7)*signed(FMAP_64_78);
			MULT_79(63)<=signed(DIN_79_7)*signed(FMAP_64_79);
			MULT_80(63)<=signed(DIN_80_7)*signed(FMAP_64_80);
			MULT_81(63)<=signed(DIN_81_7)*signed(FMAP_64_81);
			MULT_82(63)<=signed(DIN_82_7)*signed(FMAP_64_82);
			MULT_83(63)<=signed(DIN_83_7)*signed(FMAP_64_83);
			MULT_84(63)<=signed(DIN_84_7)*signed(FMAP_64_84);
			MULT_85(63)<=signed(DIN_85_7)*signed(FMAP_64_85);
			MULT_86(63)<=signed(DIN_86_7)*signed(FMAP_64_86);
			MULT_87(63)<=signed(DIN_87_7)*signed(FMAP_64_87);
			MULT_88(63)<=signed(DIN_88_7)*signed(FMAP_64_88);
			MULT_89(63)<=signed(DIN_89_7)*signed(FMAP_64_89);
			MULT_90(63)<=signed(DIN_90_7)*signed(FMAP_64_90);
			MULT_91(63)<=signed(DIN_91_7)*signed(FMAP_64_91);
			MULT_92(63)<=signed(DIN_92_7)*signed(FMAP_64_92);
			MULT_93(63)<=signed(DIN_93_7)*signed(FMAP_64_93);
			MULT_94(63)<=signed(DIN_94_7)*signed(FMAP_64_94);
			MULT_95(63)<=signed(DIN_95_7)*signed(FMAP_64_95);
			MULT_96(63)<=signed(DIN_96_7)*signed(FMAP_64_96);
			MULT_97(63)<=signed(DIN_97_7)*signed(FMAP_64_97);
			MULT_98(63)<=signed(DIN_98_7)*signed(FMAP_64_98);
			MULT_99(63)<=signed(DIN_99_7)*signed(FMAP_64_99);
			MULT_100(63)<=signed(DIN_100_7)*signed(FMAP_64_100);
			MULT_101(63)<=signed(DIN_101_7)*signed(FMAP_64_101);
			MULT_102(63)<=signed(DIN_102_7)*signed(FMAP_64_102);
			MULT_103(63)<=signed(DIN_103_7)*signed(FMAP_64_103);
			MULT_104(63)<=signed(DIN_104_7)*signed(FMAP_64_104);
			MULT_105(63)<=signed(DIN_105_7)*signed(FMAP_64_105);
			MULT_106(63)<=signed(DIN_106_7)*signed(FMAP_64_106);
			MULT_107(63)<=signed(DIN_107_7)*signed(FMAP_64_107);
			MULT_108(63)<=signed(DIN_108_7)*signed(FMAP_64_108);
			MULT_109(63)<=signed(DIN_109_7)*signed(FMAP_64_109);
			MULT_110(63)<=signed(DIN_110_7)*signed(FMAP_64_110);
			MULT_111(63)<=signed(DIN_111_7)*signed(FMAP_64_111);
			MULT_112(63)<=signed(DIN_112_7)*signed(FMAP_64_112);
			MULT_113(63)<=signed(DIN_113_7)*signed(FMAP_64_113);
			MULT_114(63)<=signed(DIN_114_7)*signed(FMAP_64_114);
			MULT_115(63)<=signed(DIN_115_7)*signed(FMAP_64_115);
			MULT_116(63)<=signed(DIN_116_7)*signed(FMAP_64_116);
			MULT_117(63)<=signed(DIN_117_7)*signed(FMAP_64_117);
			MULT_118(63)<=signed(DIN_118_7)*signed(FMAP_64_118);
			MULT_119(63)<=signed(DIN_119_7)*signed(FMAP_64_119);
			MULT_120(63)<=signed(DIN_120_7)*signed(FMAP_64_120);

			MULT_1(64)<=signed(DIN_1_7)*signed(FMAP_65_1);
			MULT_2(64)<=signed(DIN_2_7)*signed(FMAP_65_2);
			MULT_3(64)<=signed(DIN_3_7)*signed(FMAP_65_3);
			MULT_4(64)<=signed(DIN_4_7)*signed(FMAP_65_4);
			MULT_5(64)<=signed(DIN_5_7)*signed(FMAP_65_5);
			MULT_6(64)<=signed(DIN_6_7)*signed(FMAP_65_6);
			MULT_7(64)<=signed(DIN_7_7)*signed(FMAP_65_7);
			MULT_8(64)<=signed(DIN_8_7)*signed(FMAP_65_8);
			MULT_9(64)<=signed(DIN_9_7)*signed(FMAP_65_9);
			MULT_10(64)<=signed(DIN_10_7)*signed(FMAP_65_10);
			MULT_11(64)<=signed(DIN_11_7)*signed(FMAP_65_11);
			MULT_12(64)<=signed(DIN_12_7)*signed(FMAP_65_12);
			MULT_13(64)<=signed(DIN_13_7)*signed(FMAP_65_13);
			MULT_14(64)<=signed(DIN_14_7)*signed(FMAP_65_14);
			MULT_15(64)<=signed(DIN_15_7)*signed(FMAP_65_15);
			MULT_16(64)<=signed(DIN_16_7)*signed(FMAP_65_16);
			MULT_17(64)<=signed(DIN_17_7)*signed(FMAP_65_17);
			MULT_18(64)<=signed(DIN_18_7)*signed(FMAP_65_18);
			MULT_19(64)<=signed(DIN_19_7)*signed(FMAP_65_19);
			MULT_20(64)<=signed(DIN_20_7)*signed(FMAP_65_20);
			MULT_21(64)<=signed(DIN_21_7)*signed(FMAP_65_21);
			MULT_22(64)<=signed(DIN_22_7)*signed(FMAP_65_22);
			MULT_23(64)<=signed(DIN_23_7)*signed(FMAP_65_23);
			MULT_24(64)<=signed(DIN_24_7)*signed(FMAP_65_24);
			MULT_25(64)<=signed(DIN_25_7)*signed(FMAP_65_25);
			MULT_26(64)<=signed(DIN_26_7)*signed(FMAP_65_26);
			MULT_27(64)<=signed(DIN_27_7)*signed(FMAP_65_27);
			MULT_28(64)<=signed(DIN_28_7)*signed(FMAP_65_28);
			MULT_29(64)<=signed(DIN_29_7)*signed(FMAP_65_29);
			MULT_30(64)<=signed(DIN_30_7)*signed(FMAP_65_30);
			MULT_31(64)<=signed(DIN_31_7)*signed(FMAP_65_31);
			MULT_32(64)<=signed(DIN_32_7)*signed(FMAP_65_32);
			MULT_33(64)<=signed(DIN_33_7)*signed(FMAP_65_33);
			MULT_34(64)<=signed(DIN_34_7)*signed(FMAP_65_34);
			MULT_35(64)<=signed(DIN_35_7)*signed(FMAP_65_35);
			MULT_36(64)<=signed(DIN_36_7)*signed(FMAP_65_36);
			MULT_37(64)<=signed(DIN_37_7)*signed(FMAP_65_37);
			MULT_38(64)<=signed(DIN_38_7)*signed(FMAP_65_38);
			MULT_39(64)<=signed(DIN_39_7)*signed(FMAP_65_39);
			MULT_40(64)<=signed(DIN_40_7)*signed(FMAP_65_40);
			MULT_41(64)<=signed(DIN_41_7)*signed(FMAP_65_41);
			MULT_42(64)<=signed(DIN_42_7)*signed(FMAP_65_42);
			MULT_43(64)<=signed(DIN_43_7)*signed(FMAP_65_43);
			MULT_44(64)<=signed(DIN_44_7)*signed(FMAP_65_44);
			MULT_45(64)<=signed(DIN_45_7)*signed(FMAP_65_45);
			MULT_46(64)<=signed(DIN_46_7)*signed(FMAP_65_46);
			MULT_47(64)<=signed(DIN_47_7)*signed(FMAP_65_47);
			MULT_48(64)<=signed(DIN_48_7)*signed(FMAP_65_48);
			MULT_49(64)<=signed(DIN_49_7)*signed(FMAP_65_49);
			MULT_50(64)<=signed(DIN_50_7)*signed(FMAP_65_50);
			MULT_51(64)<=signed(DIN_51_7)*signed(FMAP_65_51);
			MULT_52(64)<=signed(DIN_52_7)*signed(FMAP_65_52);
			MULT_53(64)<=signed(DIN_53_7)*signed(FMAP_65_53);
			MULT_54(64)<=signed(DIN_54_7)*signed(FMAP_65_54);
			MULT_55(64)<=signed(DIN_55_7)*signed(FMAP_65_55);
			MULT_56(64)<=signed(DIN_56_7)*signed(FMAP_65_56);
			MULT_57(64)<=signed(DIN_57_7)*signed(FMAP_65_57);
			MULT_58(64)<=signed(DIN_58_7)*signed(FMAP_65_58);
			MULT_59(64)<=signed(DIN_59_7)*signed(FMAP_65_59);
			MULT_60(64)<=signed(DIN_60_7)*signed(FMAP_65_60);
			MULT_61(64)<=signed(DIN_61_7)*signed(FMAP_65_61);
			MULT_62(64)<=signed(DIN_62_7)*signed(FMAP_65_62);
			MULT_63(64)<=signed(DIN_63_7)*signed(FMAP_65_63);
			MULT_64(64)<=signed(DIN_64_7)*signed(FMAP_65_64);
			MULT_65(64)<=signed(DIN_65_7)*signed(FMAP_65_65);
			MULT_66(64)<=signed(DIN_66_7)*signed(FMAP_65_66);
			MULT_67(64)<=signed(DIN_67_7)*signed(FMAP_65_67);
			MULT_68(64)<=signed(DIN_68_7)*signed(FMAP_65_68);
			MULT_69(64)<=signed(DIN_69_7)*signed(FMAP_65_69);
			MULT_70(64)<=signed(DIN_70_7)*signed(FMAP_65_70);
			MULT_71(64)<=signed(DIN_71_7)*signed(FMAP_65_71);
			MULT_72(64)<=signed(DIN_72_7)*signed(FMAP_65_72);
			MULT_73(64)<=signed(DIN_73_7)*signed(FMAP_65_73);
			MULT_74(64)<=signed(DIN_74_7)*signed(FMAP_65_74);
			MULT_75(64)<=signed(DIN_75_7)*signed(FMAP_65_75);
			MULT_76(64)<=signed(DIN_76_7)*signed(FMAP_65_76);
			MULT_77(64)<=signed(DIN_77_7)*signed(FMAP_65_77);
			MULT_78(64)<=signed(DIN_78_7)*signed(FMAP_65_78);
			MULT_79(64)<=signed(DIN_79_7)*signed(FMAP_65_79);
			MULT_80(64)<=signed(DIN_80_7)*signed(FMAP_65_80);
			MULT_81(64)<=signed(DIN_81_7)*signed(FMAP_65_81);
			MULT_82(64)<=signed(DIN_82_7)*signed(FMAP_65_82);
			MULT_83(64)<=signed(DIN_83_7)*signed(FMAP_65_83);
			MULT_84(64)<=signed(DIN_84_7)*signed(FMAP_65_84);
			MULT_85(64)<=signed(DIN_85_7)*signed(FMAP_65_85);
			MULT_86(64)<=signed(DIN_86_7)*signed(FMAP_65_86);
			MULT_87(64)<=signed(DIN_87_7)*signed(FMAP_65_87);
			MULT_88(64)<=signed(DIN_88_7)*signed(FMAP_65_88);
			MULT_89(64)<=signed(DIN_89_7)*signed(FMAP_65_89);
			MULT_90(64)<=signed(DIN_90_7)*signed(FMAP_65_90);
			MULT_91(64)<=signed(DIN_91_7)*signed(FMAP_65_91);
			MULT_92(64)<=signed(DIN_92_7)*signed(FMAP_65_92);
			MULT_93(64)<=signed(DIN_93_7)*signed(FMAP_65_93);
			MULT_94(64)<=signed(DIN_94_7)*signed(FMAP_65_94);
			MULT_95(64)<=signed(DIN_95_7)*signed(FMAP_65_95);
			MULT_96(64)<=signed(DIN_96_7)*signed(FMAP_65_96);
			MULT_97(64)<=signed(DIN_97_7)*signed(FMAP_65_97);
			MULT_98(64)<=signed(DIN_98_7)*signed(FMAP_65_98);
			MULT_99(64)<=signed(DIN_99_7)*signed(FMAP_65_99);
			MULT_100(64)<=signed(DIN_100_7)*signed(FMAP_65_100);
			MULT_101(64)<=signed(DIN_101_7)*signed(FMAP_65_101);
			MULT_102(64)<=signed(DIN_102_7)*signed(FMAP_65_102);
			MULT_103(64)<=signed(DIN_103_7)*signed(FMAP_65_103);
			MULT_104(64)<=signed(DIN_104_7)*signed(FMAP_65_104);
			MULT_105(64)<=signed(DIN_105_7)*signed(FMAP_65_105);
			MULT_106(64)<=signed(DIN_106_7)*signed(FMAP_65_106);
			MULT_107(64)<=signed(DIN_107_7)*signed(FMAP_65_107);
			MULT_108(64)<=signed(DIN_108_7)*signed(FMAP_65_108);
			MULT_109(64)<=signed(DIN_109_7)*signed(FMAP_65_109);
			MULT_110(64)<=signed(DIN_110_7)*signed(FMAP_65_110);
			MULT_111(64)<=signed(DIN_111_7)*signed(FMAP_65_111);
			MULT_112(64)<=signed(DIN_112_7)*signed(FMAP_65_112);
			MULT_113(64)<=signed(DIN_113_7)*signed(FMAP_65_113);
			MULT_114(64)<=signed(DIN_114_7)*signed(FMAP_65_114);
			MULT_115(64)<=signed(DIN_115_7)*signed(FMAP_65_115);
			MULT_116(64)<=signed(DIN_116_7)*signed(FMAP_65_116);
			MULT_117(64)<=signed(DIN_117_7)*signed(FMAP_65_117);
			MULT_118(64)<=signed(DIN_118_7)*signed(FMAP_65_118);
			MULT_119(64)<=signed(DIN_119_7)*signed(FMAP_65_119);
			MULT_120(64)<=signed(DIN_120_7)*signed(FMAP_65_120);

			MULT_1(65)<=signed(DIN_1_7)*signed(FMAP_66_1);
			MULT_2(65)<=signed(DIN_2_7)*signed(FMAP_66_2);
			MULT_3(65)<=signed(DIN_3_7)*signed(FMAP_66_3);
			MULT_4(65)<=signed(DIN_4_7)*signed(FMAP_66_4);
			MULT_5(65)<=signed(DIN_5_7)*signed(FMAP_66_5);
			MULT_6(65)<=signed(DIN_6_7)*signed(FMAP_66_6);
			MULT_7(65)<=signed(DIN_7_7)*signed(FMAP_66_7);
			MULT_8(65)<=signed(DIN_8_7)*signed(FMAP_66_8);
			MULT_9(65)<=signed(DIN_9_7)*signed(FMAP_66_9);
			MULT_10(65)<=signed(DIN_10_7)*signed(FMAP_66_10);
			MULT_11(65)<=signed(DIN_11_7)*signed(FMAP_66_11);
			MULT_12(65)<=signed(DIN_12_7)*signed(FMAP_66_12);
			MULT_13(65)<=signed(DIN_13_7)*signed(FMAP_66_13);
			MULT_14(65)<=signed(DIN_14_7)*signed(FMAP_66_14);
			MULT_15(65)<=signed(DIN_15_7)*signed(FMAP_66_15);
			MULT_16(65)<=signed(DIN_16_7)*signed(FMAP_66_16);
			MULT_17(65)<=signed(DIN_17_7)*signed(FMAP_66_17);
			MULT_18(65)<=signed(DIN_18_7)*signed(FMAP_66_18);
			MULT_19(65)<=signed(DIN_19_7)*signed(FMAP_66_19);
			MULT_20(65)<=signed(DIN_20_7)*signed(FMAP_66_20);
			MULT_21(65)<=signed(DIN_21_7)*signed(FMAP_66_21);
			MULT_22(65)<=signed(DIN_22_7)*signed(FMAP_66_22);
			MULT_23(65)<=signed(DIN_23_7)*signed(FMAP_66_23);
			MULT_24(65)<=signed(DIN_24_7)*signed(FMAP_66_24);
			MULT_25(65)<=signed(DIN_25_7)*signed(FMAP_66_25);
			MULT_26(65)<=signed(DIN_26_7)*signed(FMAP_66_26);
			MULT_27(65)<=signed(DIN_27_7)*signed(FMAP_66_27);
			MULT_28(65)<=signed(DIN_28_7)*signed(FMAP_66_28);
			MULT_29(65)<=signed(DIN_29_7)*signed(FMAP_66_29);
			MULT_30(65)<=signed(DIN_30_7)*signed(FMAP_66_30);
			MULT_31(65)<=signed(DIN_31_7)*signed(FMAP_66_31);
			MULT_32(65)<=signed(DIN_32_7)*signed(FMAP_66_32);
			MULT_33(65)<=signed(DIN_33_7)*signed(FMAP_66_33);
			MULT_34(65)<=signed(DIN_34_7)*signed(FMAP_66_34);
			MULT_35(65)<=signed(DIN_35_7)*signed(FMAP_66_35);
			MULT_36(65)<=signed(DIN_36_7)*signed(FMAP_66_36);
			MULT_37(65)<=signed(DIN_37_7)*signed(FMAP_66_37);
			MULT_38(65)<=signed(DIN_38_7)*signed(FMAP_66_38);
			MULT_39(65)<=signed(DIN_39_7)*signed(FMAP_66_39);
			MULT_40(65)<=signed(DIN_40_7)*signed(FMAP_66_40);
			MULT_41(65)<=signed(DIN_41_7)*signed(FMAP_66_41);
			MULT_42(65)<=signed(DIN_42_7)*signed(FMAP_66_42);
			MULT_43(65)<=signed(DIN_43_7)*signed(FMAP_66_43);
			MULT_44(65)<=signed(DIN_44_7)*signed(FMAP_66_44);
			MULT_45(65)<=signed(DIN_45_7)*signed(FMAP_66_45);
			MULT_46(65)<=signed(DIN_46_7)*signed(FMAP_66_46);
			MULT_47(65)<=signed(DIN_47_7)*signed(FMAP_66_47);
			MULT_48(65)<=signed(DIN_48_7)*signed(FMAP_66_48);
			MULT_49(65)<=signed(DIN_49_7)*signed(FMAP_66_49);
			MULT_50(65)<=signed(DIN_50_7)*signed(FMAP_66_50);
			MULT_51(65)<=signed(DIN_51_7)*signed(FMAP_66_51);
			MULT_52(65)<=signed(DIN_52_7)*signed(FMAP_66_52);
			MULT_53(65)<=signed(DIN_53_7)*signed(FMAP_66_53);
			MULT_54(65)<=signed(DIN_54_7)*signed(FMAP_66_54);
			MULT_55(65)<=signed(DIN_55_7)*signed(FMAP_66_55);
			MULT_56(65)<=signed(DIN_56_7)*signed(FMAP_66_56);
			MULT_57(65)<=signed(DIN_57_7)*signed(FMAP_66_57);
			MULT_58(65)<=signed(DIN_58_7)*signed(FMAP_66_58);
			MULT_59(65)<=signed(DIN_59_7)*signed(FMAP_66_59);
			MULT_60(65)<=signed(DIN_60_7)*signed(FMAP_66_60);
			MULT_61(65)<=signed(DIN_61_7)*signed(FMAP_66_61);
			MULT_62(65)<=signed(DIN_62_7)*signed(FMAP_66_62);
			MULT_63(65)<=signed(DIN_63_7)*signed(FMAP_66_63);
			MULT_64(65)<=signed(DIN_64_7)*signed(FMAP_66_64);
			MULT_65(65)<=signed(DIN_65_7)*signed(FMAP_66_65);
			MULT_66(65)<=signed(DIN_66_7)*signed(FMAP_66_66);
			MULT_67(65)<=signed(DIN_67_7)*signed(FMAP_66_67);
			MULT_68(65)<=signed(DIN_68_7)*signed(FMAP_66_68);
			MULT_69(65)<=signed(DIN_69_7)*signed(FMAP_66_69);
			MULT_70(65)<=signed(DIN_70_7)*signed(FMAP_66_70);
			MULT_71(65)<=signed(DIN_71_7)*signed(FMAP_66_71);
			MULT_72(65)<=signed(DIN_72_7)*signed(FMAP_66_72);
			MULT_73(65)<=signed(DIN_73_7)*signed(FMAP_66_73);
			MULT_74(65)<=signed(DIN_74_7)*signed(FMAP_66_74);
			MULT_75(65)<=signed(DIN_75_7)*signed(FMAP_66_75);
			MULT_76(65)<=signed(DIN_76_7)*signed(FMAP_66_76);
			MULT_77(65)<=signed(DIN_77_7)*signed(FMAP_66_77);
			MULT_78(65)<=signed(DIN_78_7)*signed(FMAP_66_78);
			MULT_79(65)<=signed(DIN_79_7)*signed(FMAP_66_79);
			MULT_80(65)<=signed(DIN_80_7)*signed(FMAP_66_80);
			MULT_81(65)<=signed(DIN_81_7)*signed(FMAP_66_81);
			MULT_82(65)<=signed(DIN_82_7)*signed(FMAP_66_82);
			MULT_83(65)<=signed(DIN_83_7)*signed(FMAP_66_83);
			MULT_84(65)<=signed(DIN_84_7)*signed(FMAP_66_84);
			MULT_85(65)<=signed(DIN_85_7)*signed(FMAP_66_85);
			MULT_86(65)<=signed(DIN_86_7)*signed(FMAP_66_86);
			MULT_87(65)<=signed(DIN_87_7)*signed(FMAP_66_87);
			MULT_88(65)<=signed(DIN_88_7)*signed(FMAP_66_88);
			MULT_89(65)<=signed(DIN_89_7)*signed(FMAP_66_89);
			MULT_90(65)<=signed(DIN_90_7)*signed(FMAP_66_90);
			MULT_91(65)<=signed(DIN_91_7)*signed(FMAP_66_91);
			MULT_92(65)<=signed(DIN_92_7)*signed(FMAP_66_92);
			MULT_93(65)<=signed(DIN_93_7)*signed(FMAP_66_93);
			MULT_94(65)<=signed(DIN_94_7)*signed(FMAP_66_94);
			MULT_95(65)<=signed(DIN_95_7)*signed(FMAP_66_95);
			MULT_96(65)<=signed(DIN_96_7)*signed(FMAP_66_96);
			MULT_97(65)<=signed(DIN_97_7)*signed(FMAP_66_97);
			MULT_98(65)<=signed(DIN_98_7)*signed(FMAP_66_98);
			MULT_99(65)<=signed(DIN_99_7)*signed(FMAP_66_99);
			MULT_100(65)<=signed(DIN_100_7)*signed(FMAP_66_100);
			MULT_101(65)<=signed(DIN_101_7)*signed(FMAP_66_101);
			MULT_102(65)<=signed(DIN_102_7)*signed(FMAP_66_102);
			MULT_103(65)<=signed(DIN_103_7)*signed(FMAP_66_103);
			MULT_104(65)<=signed(DIN_104_7)*signed(FMAP_66_104);
			MULT_105(65)<=signed(DIN_105_7)*signed(FMAP_66_105);
			MULT_106(65)<=signed(DIN_106_7)*signed(FMAP_66_106);
			MULT_107(65)<=signed(DIN_107_7)*signed(FMAP_66_107);
			MULT_108(65)<=signed(DIN_108_7)*signed(FMAP_66_108);
			MULT_109(65)<=signed(DIN_109_7)*signed(FMAP_66_109);
			MULT_110(65)<=signed(DIN_110_7)*signed(FMAP_66_110);
			MULT_111(65)<=signed(DIN_111_7)*signed(FMAP_66_111);
			MULT_112(65)<=signed(DIN_112_7)*signed(FMAP_66_112);
			MULT_113(65)<=signed(DIN_113_7)*signed(FMAP_66_113);
			MULT_114(65)<=signed(DIN_114_7)*signed(FMAP_66_114);
			MULT_115(65)<=signed(DIN_115_7)*signed(FMAP_66_115);
			MULT_116(65)<=signed(DIN_116_7)*signed(FMAP_66_116);
			MULT_117(65)<=signed(DIN_117_7)*signed(FMAP_66_117);
			MULT_118(65)<=signed(DIN_118_7)*signed(FMAP_66_118);
			MULT_119(65)<=signed(DIN_119_7)*signed(FMAP_66_119);
			MULT_120(65)<=signed(DIN_120_7)*signed(FMAP_66_120);

			MULT_1(66)<=signed(DIN_1_7)*signed(FMAP_67_1);
			MULT_2(66)<=signed(DIN_2_7)*signed(FMAP_67_2);
			MULT_3(66)<=signed(DIN_3_7)*signed(FMAP_67_3);
			MULT_4(66)<=signed(DIN_4_7)*signed(FMAP_67_4);
			MULT_5(66)<=signed(DIN_5_7)*signed(FMAP_67_5);
			MULT_6(66)<=signed(DIN_6_7)*signed(FMAP_67_6);
			MULT_7(66)<=signed(DIN_7_7)*signed(FMAP_67_7);
			MULT_8(66)<=signed(DIN_8_7)*signed(FMAP_67_8);
			MULT_9(66)<=signed(DIN_9_7)*signed(FMAP_67_9);
			MULT_10(66)<=signed(DIN_10_7)*signed(FMAP_67_10);
			MULT_11(66)<=signed(DIN_11_7)*signed(FMAP_67_11);
			MULT_12(66)<=signed(DIN_12_7)*signed(FMAP_67_12);
			MULT_13(66)<=signed(DIN_13_7)*signed(FMAP_67_13);
			MULT_14(66)<=signed(DIN_14_7)*signed(FMAP_67_14);
			MULT_15(66)<=signed(DIN_15_7)*signed(FMAP_67_15);
			MULT_16(66)<=signed(DIN_16_7)*signed(FMAP_67_16);
			MULT_17(66)<=signed(DIN_17_7)*signed(FMAP_67_17);
			MULT_18(66)<=signed(DIN_18_7)*signed(FMAP_67_18);
			MULT_19(66)<=signed(DIN_19_7)*signed(FMAP_67_19);
			MULT_20(66)<=signed(DIN_20_7)*signed(FMAP_67_20);
			MULT_21(66)<=signed(DIN_21_7)*signed(FMAP_67_21);
			MULT_22(66)<=signed(DIN_22_7)*signed(FMAP_67_22);
			MULT_23(66)<=signed(DIN_23_7)*signed(FMAP_67_23);
			MULT_24(66)<=signed(DIN_24_7)*signed(FMAP_67_24);
			MULT_25(66)<=signed(DIN_25_7)*signed(FMAP_67_25);
			MULT_26(66)<=signed(DIN_26_7)*signed(FMAP_67_26);
			MULT_27(66)<=signed(DIN_27_7)*signed(FMAP_67_27);
			MULT_28(66)<=signed(DIN_28_7)*signed(FMAP_67_28);
			MULT_29(66)<=signed(DIN_29_7)*signed(FMAP_67_29);
			MULT_30(66)<=signed(DIN_30_7)*signed(FMAP_67_30);
			MULT_31(66)<=signed(DIN_31_7)*signed(FMAP_67_31);
			MULT_32(66)<=signed(DIN_32_7)*signed(FMAP_67_32);
			MULT_33(66)<=signed(DIN_33_7)*signed(FMAP_67_33);
			MULT_34(66)<=signed(DIN_34_7)*signed(FMAP_67_34);
			MULT_35(66)<=signed(DIN_35_7)*signed(FMAP_67_35);
			MULT_36(66)<=signed(DIN_36_7)*signed(FMAP_67_36);
			MULT_37(66)<=signed(DIN_37_7)*signed(FMAP_67_37);
			MULT_38(66)<=signed(DIN_38_7)*signed(FMAP_67_38);
			MULT_39(66)<=signed(DIN_39_7)*signed(FMAP_67_39);
			MULT_40(66)<=signed(DIN_40_7)*signed(FMAP_67_40);
			MULT_41(66)<=signed(DIN_41_7)*signed(FMAP_67_41);
			MULT_42(66)<=signed(DIN_42_7)*signed(FMAP_67_42);
			MULT_43(66)<=signed(DIN_43_7)*signed(FMAP_67_43);
			MULT_44(66)<=signed(DIN_44_7)*signed(FMAP_67_44);
			MULT_45(66)<=signed(DIN_45_7)*signed(FMAP_67_45);
			MULT_46(66)<=signed(DIN_46_7)*signed(FMAP_67_46);
			MULT_47(66)<=signed(DIN_47_7)*signed(FMAP_67_47);
			MULT_48(66)<=signed(DIN_48_7)*signed(FMAP_67_48);
			MULT_49(66)<=signed(DIN_49_7)*signed(FMAP_67_49);
			MULT_50(66)<=signed(DIN_50_7)*signed(FMAP_67_50);
			MULT_51(66)<=signed(DIN_51_7)*signed(FMAP_67_51);
			MULT_52(66)<=signed(DIN_52_7)*signed(FMAP_67_52);
			MULT_53(66)<=signed(DIN_53_7)*signed(FMAP_67_53);
			MULT_54(66)<=signed(DIN_54_7)*signed(FMAP_67_54);
			MULT_55(66)<=signed(DIN_55_7)*signed(FMAP_67_55);
			MULT_56(66)<=signed(DIN_56_7)*signed(FMAP_67_56);
			MULT_57(66)<=signed(DIN_57_7)*signed(FMAP_67_57);
			MULT_58(66)<=signed(DIN_58_7)*signed(FMAP_67_58);
			MULT_59(66)<=signed(DIN_59_7)*signed(FMAP_67_59);
			MULT_60(66)<=signed(DIN_60_7)*signed(FMAP_67_60);
			MULT_61(66)<=signed(DIN_61_7)*signed(FMAP_67_61);
			MULT_62(66)<=signed(DIN_62_7)*signed(FMAP_67_62);
			MULT_63(66)<=signed(DIN_63_7)*signed(FMAP_67_63);
			MULT_64(66)<=signed(DIN_64_7)*signed(FMAP_67_64);
			MULT_65(66)<=signed(DIN_65_7)*signed(FMAP_67_65);
			MULT_66(66)<=signed(DIN_66_7)*signed(FMAP_67_66);
			MULT_67(66)<=signed(DIN_67_7)*signed(FMAP_67_67);
			MULT_68(66)<=signed(DIN_68_7)*signed(FMAP_67_68);
			MULT_69(66)<=signed(DIN_69_7)*signed(FMAP_67_69);
			MULT_70(66)<=signed(DIN_70_7)*signed(FMAP_67_70);
			MULT_71(66)<=signed(DIN_71_7)*signed(FMAP_67_71);
			MULT_72(66)<=signed(DIN_72_7)*signed(FMAP_67_72);
			MULT_73(66)<=signed(DIN_73_7)*signed(FMAP_67_73);
			MULT_74(66)<=signed(DIN_74_7)*signed(FMAP_67_74);
			MULT_75(66)<=signed(DIN_75_7)*signed(FMAP_67_75);
			MULT_76(66)<=signed(DIN_76_7)*signed(FMAP_67_76);
			MULT_77(66)<=signed(DIN_77_7)*signed(FMAP_67_77);
			MULT_78(66)<=signed(DIN_78_7)*signed(FMAP_67_78);
			MULT_79(66)<=signed(DIN_79_7)*signed(FMAP_67_79);
			MULT_80(66)<=signed(DIN_80_7)*signed(FMAP_67_80);
			MULT_81(66)<=signed(DIN_81_7)*signed(FMAP_67_81);
			MULT_82(66)<=signed(DIN_82_7)*signed(FMAP_67_82);
			MULT_83(66)<=signed(DIN_83_7)*signed(FMAP_67_83);
			MULT_84(66)<=signed(DIN_84_7)*signed(FMAP_67_84);
			MULT_85(66)<=signed(DIN_85_7)*signed(FMAP_67_85);
			MULT_86(66)<=signed(DIN_86_7)*signed(FMAP_67_86);
			MULT_87(66)<=signed(DIN_87_7)*signed(FMAP_67_87);
			MULT_88(66)<=signed(DIN_88_7)*signed(FMAP_67_88);
			MULT_89(66)<=signed(DIN_89_7)*signed(FMAP_67_89);
			MULT_90(66)<=signed(DIN_90_7)*signed(FMAP_67_90);
			MULT_91(66)<=signed(DIN_91_7)*signed(FMAP_67_91);
			MULT_92(66)<=signed(DIN_92_7)*signed(FMAP_67_92);
			MULT_93(66)<=signed(DIN_93_7)*signed(FMAP_67_93);
			MULT_94(66)<=signed(DIN_94_7)*signed(FMAP_67_94);
			MULT_95(66)<=signed(DIN_95_7)*signed(FMAP_67_95);
			MULT_96(66)<=signed(DIN_96_7)*signed(FMAP_67_96);
			MULT_97(66)<=signed(DIN_97_7)*signed(FMAP_67_97);
			MULT_98(66)<=signed(DIN_98_7)*signed(FMAP_67_98);
			MULT_99(66)<=signed(DIN_99_7)*signed(FMAP_67_99);
			MULT_100(66)<=signed(DIN_100_7)*signed(FMAP_67_100);
			MULT_101(66)<=signed(DIN_101_7)*signed(FMAP_67_101);
			MULT_102(66)<=signed(DIN_102_7)*signed(FMAP_67_102);
			MULT_103(66)<=signed(DIN_103_7)*signed(FMAP_67_103);
			MULT_104(66)<=signed(DIN_104_7)*signed(FMAP_67_104);
			MULT_105(66)<=signed(DIN_105_7)*signed(FMAP_67_105);
			MULT_106(66)<=signed(DIN_106_7)*signed(FMAP_67_106);
			MULT_107(66)<=signed(DIN_107_7)*signed(FMAP_67_107);
			MULT_108(66)<=signed(DIN_108_7)*signed(FMAP_67_108);
			MULT_109(66)<=signed(DIN_109_7)*signed(FMAP_67_109);
			MULT_110(66)<=signed(DIN_110_7)*signed(FMAP_67_110);
			MULT_111(66)<=signed(DIN_111_7)*signed(FMAP_67_111);
			MULT_112(66)<=signed(DIN_112_7)*signed(FMAP_67_112);
			MULT_113(66)<=signed(DIN_113_7)*signed(FMAP_67_113);
			MULT_114(66)<=signed(DIN_114_7)*signed(FMAP_67_114);
			MULT_115(66)<=signed(DIN_115_7)*signed(FMAP_67_115);
			MULT_116(66)<=signed(DIN_116_7)*signed(FMAP_67_116);
			MULT_117(66)<=signed(DIN_117_7)*signed(FMAP_67_117);
			MULT_118(66)<=signed(DIN_118_7)*signed(FMAP_67_118);
			MULT_119(66)<=signed(DIN_119_7)*signed(FMAP_67_119);
			MULT_120(66)<=signed(DIN_120_7)*signed(FMAP_67_120);

			MULT_1(67)<=signed(DIN_1_7)*signed(FMAP_68_1);
			MULT_2(67)<=signed(DIN_2_7)*signed(FMAP_68_2);
			MULT_3(67)<=signed(DIN_3_7)*signed(FMAP_68_3);
			MULT_4(67)<=signed(DIN_4_7)*signed(FMAP_68_4);
			MULT_5(67)<=signed(DIN_5_7)*signed(FMAP_68_5);
			MULT_6(67)<=signed(DIN_6_7)*signed(FMAP_68_6);
			MULT_7(67)<=signed(DIN_7_7)*signed(FMAP_68_7);
			MULT_8(67)<=signed(DIN_8_7)*signed(FMAP_68_8);
			MULT_9(67)<=signed(DIN_9_7)*signed(FMAP_68_9);
			MULT_10(67)<=signed(DIN_10_7)*signed(FMAP_68_10);
			MULT_11(67)<=signed(DIN_11_7)*signed(FMAP_68_11);
			MULT_12(67)<=signed(DIN_12_7)*signed(FMAP_68_12);
			MULT_13(67)<=signed(DIN_13_7)*signed(FMAP_68_13);
			MULT_14(67)<=signed(DIN_14_7)*signed(FMAP_68_14);
			MULT_15(67)<=signed(DIN_15_7)*signed(FMAP_68_15);
			MULT_16(67)<=signed(DIN_16_7)*signed(FMAP_68_16);
			MULT_17(67)<=signed(DIN_17_7)*signed(FMAP_68_17);
			MULT_18(67)<=signed(DIN_18_7)*signed(FMAP_68_18);
			MULT_19(67)<=signed(DIN_19_7)*signed(FMAP_68_19);
			MULT_20(67)<=signed(DIN_20_7)*signed(FMAP_68_20);
			MULT_21(67)<=signed(DIN_21_7)*signed(FMAP_68_21);
			MULT_22(67)<=signed(DIN_22_7)*signed(FMAP_68_22);
			MULT_23(67)<=signed(DIN_23_7)*signed(FMAP_68_23);
			MULT_24(67)<=signed(DIN_24_7)*signed(FMAP_68_24);
			MULT_25(67)<=signed(DIN_25_7)*signed(FMAP_68_25);
			MULT_26(67)<=signed(DIN_26_7)*signed(FMAP_68_26);
			MULT_27(67)<=signed(DIN_27_7)*signed(FMAP_68_27);
			MULT_28(67)<=signed(DIN_28_7)*signed(FMAP_68_28);
			MULT_29(67)<=signed(DIN_29_7)*signed(FMAP_68_29);
			MULT_30(67)<=signed(DIN_30_7)*signed(FMAP_68_30);
			MULT_31(67)<=signed(DIN_31_7)*signed(FMAP_68_31);
			MULT_32(67)<=signed(DIN_32_7)*signed(FMAP_68_32);
			MULT_33(67)<=signed(DIN_33_7)*signed(FMAP_68_33);
			MULT_34(67)<=signed(DIN_34_7)*signed(FMAP_68_34);
			MULT_35(67)<=signed(DIN_35_7)*signed(FMAP_68_35);
			MULT_36(67)<=signed(DIN_36_7)*signed(FMAP_68_36);
			MULT_37(67)<=signed(DIN_37_7)*signed(FMAP_68_37);
			MULT_38(67)<=signed(DIN_38_7)*signed(FMAP_68_38);
			MULT_39(67)<=signed(DIN_39_7)*signed(FMAP_68_39);
			MULT_40(67)<=signed(DIN_40_7)*signed(FMAP_68_40);
			MULT_41(67)<=signed(DIN_41_7)*signed(FMAP_68_41);
			MULT_42(67)<=signed(DIN_42_7)*signed(FMAP_68_42);
			MULT_43(67)<=signed(DIN_43_7)*signed(FMAP_68_43);
			MULT_44(67)<=signed(DIN_44_7)*signed(FMAP_68_44);
			MULT_45(67)<=signed(DIN_45_7)*signed(FMAP_68_45);
			MULT_46(67)<=signed(DIN_46_7)*signed(FMAP_68_46);
			MULT_47(67)<=signed(DIN_47_7)*signed(FMAP_68_47);
			MULT_48(67)<=signed(DIN_48_7)*signed(FMAP_68_48);
			MULT_49(67)<=signed(DIN_49_7)*signed(FMAP_68_49);
			MULT_50(67)<=signed(DIN_50_7)*signed(FMAP_68_50);
			MULT_51(67)<=signed(DIN_51_7)*signed(FMAP_68_51);
			MULT_52(67)<=signed(DIN_52_7)*signed(FMAP_68_52);
			MULT_53(67)<=signed(DIN_53_7)*signed(FMAP_68_53);
			MULT_54(67)<=signed(DIN_54_7)*signed(FMAP_68_54);
			MULT_55(67)<=signed(DIN_55_7)*signed(FMAP_68_55);
			MULT_56(67)<=signed(DIN_56_7)*signed(FMAP_68_56);
			MULT_57(67)<=signed(DIN_57_7)*signed(FMAP_68_57);
			MULT_58(67)<=signed(DIN_58_7)*signed(FMAP_68_58);
			MULT_59(67)<=signed(DIN_59_7)*signed(FMAP_68_59);
			MULT_60(67)<=signed(DIN_60_7)*signed(FMAP_68_60);
			MULT_61(67)<=signed(DIN_61_7)*signed(FMAP_68_61);
			MULT_62(67)<=signed(DIN_62_7)*signed(FMAP_68_62);
			MULT_63(67)<=signed(DIN_63_7)*signed(FMAP_68_63);
			MULT_64(67)<=signed(DIN_64_7)*signed(FMAP_68_64);
			MULT_65(67)<=signed(DIN_65_7)*signed(FMAP_68_65);
			MULT_66(67)<=signed(DIN_66_7)*signed(FMAP_68_66);
			MULT_67(67)<=signed(DIN_67_7)*signed(FMAP_68_67);
			MULT_68(67)<=signed(DIN_68_7)*signed(FMAP_68_68);
			MULT_69(67)<=signed(DIN_69_7)*signed(FMAP_68_69);
			MULT_70(67)<=signed(DIN_70_7)*signed(FMAP_68_70);
			MULT_71(67)<=signed(DIN_71_7)*signed(FMAP_68_71);
			MULT_72(67)<=signed(DIN_72_7)*signed(FMAP_68_72);
			MULT_73(67)<=signed(DIN_73_7)*signed(FMAP_68_73);
			MULT_74(67)<=signed(DIN_74_7)*signed(FMAP_68_74);
			MULT_75(67)<=signed(DIN_75_7)*signed(FMAP_68_75);
			MULT_76(67)<=signed(DIN_76_7)*signed(FMAP_68_76);
			MULT_77(67)<=signed(DIN_77_7)*signed(FMAP_68_77);
			MULT_78(67)<=signed(DIN_78_7)*signed(FMAP_68_78);
			MULT_79(67)<=signed(DIN_79_7)*signed(FMAP_68_79);
			MULT_80(67)<=signed(DIN_80_7)*signed(FMAP_68_80);
			MULT_81(67)<=signed(DIN_81_7)*signed(FMAP_68_81);
			MULT_82(67)<=signed(DIN_82_7)*signed(FMAP_68_82);
			MULT_83(67)<=signed(DIN_83_7)*signed(FMAP_68_83);
			MULT_84(67)<=signed(DIN_84_7)*signed(FMAP_68_84);
			MULT_85(67)<=signed(DIN_85_7)*signed(FMAP_68_85);
			MULT_86(67)<=signed(DIN_86_7)*signed(FMAP_68_86);
			MULT_87(67)<=signed(DIN_87_7)*signed(FMAP_68_87);
			MULT_88(67)<=signed(DIN_88_7)*signed(FMAP_68_88);
			MULT_89(67)<=signed(DIN_89_7)*signed(FMAP_68_89);
			MULT_90(67)<=signed(DIN_90_7)*signed(FMAP_68_90);
			MULT_91(67)<=signed(DIN_91_7)*signed(FMAP_68_91);
			MULT_92(67)<=signed(DIN_92_7)*signed(FMAP_68_92);
			MULT_93(67)<=signed(DIN_93_7)*signed(FMAP_68_93);
			MULT_94(67)<=signed(DIN_94_7)*signed(FMAP_68_94);
			MULT_95(67)<=signed(DIN_95_7)*signed(FMAP_68_95);
			MULT_96(67)<=signed(DIN_96_7)*signed(FMAP_68_96);
			MULT_97(67)<=signed(DIN_97_7)*signed(FMAP_68_97);
			MULT_98(67)<=signed(DIN_98_7)*signed(FMAP_68_98);
			MULT_99(67)<=signed(DIN_99_7)*signed(FMAP_68_99);
			MULT_100(67)<=signed(DIN_100_7)*signed(FMAP_68_100);
			MULT_101(67)<=signed(DIN_101_7)*signed(FMAP_68_101);
			MULT_102(67)<=signed(DIN_102_7)*signed(FMAP_68_102);
			MULT_103(67)<=signed(DIN_103_7)*signed(FMAP_68_103);
			MULT_104(67)<=signed(DIN_104_7)*signed(FMAP_68_104);
			MULT_105(67)<=signed(DIN_105_7)*signed(FMAP_68_105);
			MULT_106(67)<=signed(DIN_106_7)*signed(FMAP_68_106);
			MULT_107(67)<=signed(DIN_107_7)*signed(FMAP_68_107);
			MULT_108(67)<=signed(DIN_108_7)*signed(FMAP_68_108);
			MULT_109(67)<=signed(DIN_109_7)*signed(FMAP_68_109);
			MULT_110(67)<=signed(DIN_110_7)*signed(FMAP_68_110);
			MULT_111(67)<=signed(DIN_111_7)*signed(FMAP_68_111);
			MULT_112(67)<=signed(DIN_112_7)*signed(FMAP_68_112);
			MULT_113(67)<=signed(DIN_113_7)*signed(FMAP_68_113);
			MULT_114(67)<=signed(DIN_114_7)*signed(FMAP_68_114);
			MULT_115(67)<=signed(DIN_115_7)*signed(FMAP_68_115);
			MULT_116(67)<=signed(DIN_116_7)*signed(FMAP_68_116);
			MULT_117(67)<=signed(DIN_117_7)*signed(FMAP_68_117);
			MULT_118(67)<=signed(DIN_118_7)*signed(FMAP_68_118);
			MULT_119(67)<=signed(DIN_119_7)*signed(FMAP_68_119);
			MULT_120(67)<=signed(DIN_120_7)*signed(FMAP_68_120);

			MULT_1(68)<=signed(DIN_1_7)*signed(FMAP_69_1);
			MULT_2(68)<=signed(DIN_2_7)*signed(FMAP_69_2);
			MULT_3(68)<=signed(DIN_3_7)*signed(FMAP_69_3);
			MULT_4(68)<=signed(DIN_4_7)*signed(FMAP_69_4);
			MULT_5(68)<=signed(DIN_5_7)*signed(FMAP_69_5);
			MULT_6(68)<=signed(DIN_6_7)*signed(FMAP_69_6);
			MULT_7(68)<=signed(DIN_7_7)*signed(FMAP_69_7);
			MULT_8(68)<=signed(DIN_8_7)*signed(FMAP_69_8);
			MULT_9(68)<=signed(DIN_9_7)*signed(FMAP_69_9);
			MULT_10(68)<=signed(DIN_10_7)*signed(FMAP_69_10);
			MULT_11(68)<=signed(DIN_11_7)*signed(FMAP_69_11);
			MULT_12(68)<=signed(DIN_12_7)*signed(FMAP_69_12);
			MULT_13(68)<=signed(DIN_13_7)*signed(FMAP_69_13);
			MULT_14(68)<=signed(DIN_14_7)*signed(FMAP_69_14);
			MULT_15(68)<=signed(DIN_15_7)*signed(FMAP_69_15);
			MULT_16(68)<=signed(DIN_16_7)*signed(FMAP_69_16);
			MULT_17(68)<=signed(DIN_17_7)*signed(FMAP_69_17);
			MULT_18(68)<=signed(DIN_18_7)*signed(FMAP_69_18);
			MULT_19(68)<=signed(DIN_19_7)*signed(FMAP_69_19);
			MULT_20(68)<=signed(DIN_20_7)*signed(FMAP_69_20);
			MULT_21(68)<=signed(DIN_21_7)*signed(FMAP_69_21);
			MULT_22(68)<=signed(DIN_22_7)*signed(FMAP_69_22);
			MULT_23(68)<=signed(DIN_23_7)*signed(FMAP_69_23);
			MULT_24(68)<=signed(DIN_24_7)*signed(FMAP_69_24);
			MULT_25(68)<=signed(DIN_25_7)*signed(FMAP_69_25);
			MULT_26(68)<=signed(DIN_26_7)*signed(FMAP_69_26);
			MULT_27(68)<=signed(DIN_27_7)*signed(FMAP_69_27);
			MULT_28(68)<=signed(DIN_28_7)*signed(FMAP_69_28);
			MULT_29(68)<=signed(DIN_29_7)*signed(FMAP_69_29);
			MULT_30(68)<=signed(DIN_30_7)*signed(FMAP_69_30);
			MULT_31(68)<=signed(DIN_31_7)*signed(FMAP_69_31);
			MULT_32(68)<=signed(DIN_32_7)*signed(FMAP_69_32);
			MULT_33(68)<=signed(DIN_33_7)*signed(FMAP_69_33);
			MULT_34(68)<=signed(DIN_34_7)*signed(FMAP_69_34);
			MULT_35(68)<=signed(DIN_35_7)*signed(FMAP_69_35);
			MULT_36(68)<=signed(DIN_36_7)*signed(FMAP_69_36);
			MULT_37(68)<=signed(DIN_37_7)*signed(FMAP_69_37);
			MULT_38(68)<=signed(DIN_38_7)*signed(FMAP_69_38);
			MULT_39(68)<=signed(DIN_39_7)*signed(FMAP_69_39);
			MULT_40(68)<=signed(DIN_40_7)*signed(FMAP_69_40);
			MULT_41(68)<=signed(DIN_41_7)*signed(FMAP_69_41);
			MULT_42(68)<=signed(DIN_42_7)*signed(FMAP_69_42);
			MULT_43(68)<=signed(DIN_43_7)*signed(FMAP_69_43);
			MULT_44(68)<=signed(DIN_44_7)*signed(FMAP_69_44);
			MULT_45(68)<=signed(DIN_45_7)*signed(FMAP_69_45);
			MULT_46(68)<=signed(DIN_46_7)*signed(FMAP_69_46);
			MULT_47(68)<=signed(DIN_47_7)*signed(FMAP_69_47);
			MULT_48(68)<=signed(DIN_48_7)*signed(FMAP_69_48);
			MULT_49(68)<=signed(DIN_49_7)*signed(FMAP_69_49);
			MULT_50(68)<=signed(DIN_50_7)*signed(FMAP_69_50);
			MULT_51(68)<=signed(DIN_51_7)*signed(FMAP_69_51);
			MULT_52(68)<=signed(DIN_52_7)*signed(FMAP_69_52);
			MULT_53(68)<=signed(DIN_53_7)*signed(FMAP_69_53);
			MULT_54(68)<=signed(DIN_54_7)*signed(FMAP_69_54);
			MULT_55(68)<=signed(DIN_55_7)*signed(FMAP_69_55);
			MULT_56(68)<=signed(DIN_56_7)*signed(FMAP_69_56);
			MULT_57(68)<=signed(DIN_57_7)*signed(FMAP_69_57);
			MULT_58(68)<=signed(DIN_58_7)*signed(FMAP_69_58);
			MULT_59(68)<=signed(DIN_59_7)*signed(FMAP_69_59);
			MULT_60(68)<=signed(DIN_60_7)*signed(FMAP_69_60);
			MULT_61(68)<=signed(DIN_61_7)*signed(FMAP_69_61);
			MULT_62(68)<=signed(DIN_62_7)*signed(FMAP_69_62);
			MULT_63(68)<=signed(DIN_63_7)*signed(FMAP_69_63);
			MULT_64(68)<=signed(DIN_64_7)*signed(FMAP_69_64);
			MULT_65(68)<=signed(DIN_65_7)*signed(FMAP_69_65);
			MULT_66(68)<=signed(DIN_66_7)*signed(FMAP_69_66);
			MULT_67(68)<=signed(DIN_67_7)*signed(FMAP_69_67);
			MULT_68(68)<=signed(DIN_68_7)*signed(FMAP_69_68);
			MULT_69(68)<=signed(DIN_69_7)*signed(FMAP_69_69);
			MULT_70(68)<=signed(DIN_70_7)*signed(FMAP_69_70);
			MULT_71(68)<=signed(DIN_71_7)*signed(FMAP_69_71);
			MULT_72(68)<=signed(DIN_72_7)*signed(FMAP_69_72);
			MULT_73(68)<=signed(DIN_73_7)*signed(FMAP_69_73);
			MULT_74(68)<=signed(DIN_74_7)*signed(FMAP_69_74);
			MULT_75(68)<=signed(DIN_75_7)*signed(FMAP_69_75);
			MULT_76(68)<=signed(DIN_76_7)*signed(FMAP_69_76);
			MULT_77(68)<=signed(DIN_77_7)*signed(FMAP_69_77);
			MULT_78(68)<=signed(DIN_78_7)*signed(FMAP_69_78);
			MULT_79(68)<=signed(DIN_79_7)*signed(FMAP_69_79);
			MULT_80(68)<=signed(DIN_80_7)*signed(FMAP_69_80);
			MULT_81(68)<=signed(DIN_81_7)*signed(FMAP_69_81);
			MULT_82(68)<=signed(DIN_82_7)*signed(FMAP_69_82);
			MULT_83(68)<=signed(DIN_83_7)*signed(FMAP_69_83);
			MULT_84(68)<=signed(DIN_84_7)*signed(FMAP_69_84);
			MULT_85(68)<=signed(DIN_85_7)*signed(FMAP_69_85);
			MULT_86(68)<=signed(DIN_86_7)*signed(FMAP_69_86);
			MULT_87(68)<=signed(DIN_87_7)*signed(FMAP_69_87);
			MULT_88(68)<=signed(DIN_88_7)*signed(FMAP_69_88);
			MULT_89(68)<=signed(DIN_89_7)*signed(FMAP_69_89);
			MULT_90(68)<=signed(DIN_90_7)*signed(FMAP_69_90);
			MULT_91(68)<=signed(DIN_91_7)*signed(FMAP_69_91);
			MULT_92(68)<=signed(DIN_92_7)*signed(FMAP_69_92);
			MULT_93(68)<=signed(DIN_93_7)*signed(FMAP_69_93);
			MULT_94(68)<=signed(DIN_94_7)*signed(FMAP_69_94);
			MULT_95(68)<=signed(DIN_95_7)*signed(FMAP_69_95);
			MULT_96(68)<=signed(DIN_96_7)*signed(FMAP_69_96);
			MULT_97(68)<=signed(DIN_97_7)*signed(FMAP_69_97);
			MULT_98(68)<=signed(DIN_98_7)*signed(FMAP_69_98);
			MULT_99(68)<=signed(DIN_99_7)*signed(FMAP_69_99);
			MULT_100(68)<=signed(DIN_100_7)*signed(FMAP_69_100);
			MULT_101(68)<=signed(DIN_101_7)*signed(FMAP_69_101);
			MULT_102(68)<=signed(DIN_102_7)*signed(FMAP_69_102);
			MULT_103(68)<=signed(DIN_103_7)*signed(FMAP_69_103);
			MULT_104(68)<=signed(DIN_104_7)*signed(FMAP_69_104);
			MULT_105(68)<=signed(DIN_105_7)*signed(FMAP_69_105);
			MULT_106(68)<=signed(DIN_106_7)*signed(FMAP_69_106);
			MULT_107(68)<=signed(DIN_107_7)*signed(FMAP_69_107);
			MULT_108(68)<=signed(DIN_108_7)*signed(FMAP_69_108);
			MULT_109(68)<=signed(DIN_109_7)*signed(FMAP_69_109);
			MULT_110(68)<=signed(DIN_110_7)*signed(FMAP_69_110);
			MULT_111(68)<=signed(DIN_111_7)*signed(FMAP_69_111);
			MULT_112(68)<=signed(DIN_112_7)*signed(FMAP_69_112);
			MULT_113(68)<=signed(DIN_113_7)*signed(FMAP_69_113);
			MULT_114(68)<=signed(DIN_114_7)*signed(FMAP_69_114);
			MULT_115(68)<=signed(DIN_115_7)*signed(FMAP_69_115);
			MULT_116(68)<=signed(DIN_116_7)*signed(FMAP_69_116);
			MULT_117(68)<=signed(DIN_117_7)*signed(FMAP_69_117);
			MULT_118(68)<=signed(DIN_118_7)*signed(FMAP_69_118);
			MULT_119(68)<=signed(DIN_119_7)*signed(FMAP_69_119);
			MULT_120(68)<=signed(DIN_120_7)*signed(FMAP_69_120);

			MULT_1(69)<=signed(DIN_1_7)*signed(FMAP_70_1);
			MULT_2(69)<=signed(DIN_2_7)*signed(FMAP_70_2);
			MULT_3(69)<=signed(DIN_3_7)*signed(FMAP_70_3);
			MULT_4(69)<=signed(DIN_4_7)*signed(FMAP_70_4);
			MULT_5(69)<=signed(DIN_5_7)*signed(FMAP_70_5);
			MULT_6(69)<=signed(DIN_6_7)*signed(FMAP_70_6);
			MULT_7(69)<=signed(DIN_7_7)*signed(FMAP_70_7);
			MULT_8(69)<=signed(DIN_8_7)*signed(FMAP_70_8);
			MULT_9(69)<=signed(DIN_9_7)*signed(FMAP_70_9);
			MULT_10(69)<=signed(DIN_10_7)*signed(FMAP_70_10);
			MULT_11(69)<=signed(DIN_11_7)*signed(FMAP_70_11);
			MULT_12(69)<=signed(DIN_12_7)*signed(FMAP_70_12);
			MULT_13(69)<=signed(DIN_13_7)*signed(FMAP_70_13);
			MULT_14(69)<=signed(DIN_14_7)*signed(FMAP_70_14);
			MULT_15(69)<=signed(DIN_15_7)*signed(FMAP_70_15);
			MULT_16(69)<=signed(DIN_16_7)*signed(FMAP_70_16);
			MULT_17(69)<=signed(DIN_17_7)*signed(FMAP_70_17);
			MULT_18(69)<=signed(DIN_18_7)*signed(FMAP_70_18);
			MULT_19(69)<=signed(DIN_19_7)*signed(FMAP_70_19);
			MULT_20(69)<=signed(DIN_20_7)*signed(FMAP_70_20);
			MULT_21(69)<=signed(DIN_21_7)*signed(FMAP_70_21);
			MULT_22(69)<=signed(DIN_22_7)*signed(FMAP_70_22);
			MULT_23(69)<=signed(DIN_23_7)*signed(FMAP_70_23);
			MULT_24(69)<=signed(DIN_24_7)*signed(FMAP_70_24);
			MULT_25(69)<=signed(DIN_25_7)*signed(FMAP_70_25);
			MULT_26(69)<=signed(DIN_26_7)*signed(FMAP_70_26);
			MULT_27(69)<=signed(DIN_27_7)*signed(FMAP_70_27);
			MULT_28(69)<=signed(DIN_28_7)*signed(FMAP_70_28);
			MULT_29(69)<=signed(DIN_29_7)*signed(FMAP_70_29);
			MULT_30(69)<=signed(DIN_30_7)*signed(FMAP_70_30);
			MULT_31(69)<=signed(DIN_31_7)*signed(FMAP_70_31);
			MULT_32(69)<=signed(DIN_32_7)*signed(FMAP_70_32);
			MULT_33(69)<=signed(DIN_33_7)*signed(FMAP_70_33);
			MULT_34(69)<=signed(DIN_34_7)*signed(FMAP_70_34);
			MULT_35(69)<=signed(DIN_35_7)*signed(FMAP_70_35);
			MULT_36(69)<=signed(DIN_36_7)*signed(FMAP_70_36);
			MULT_37(69)<=signed(DIN_37_7)*signed(FMAP_70_37);
			MULT_38(69)<=signed(DIN_38_7)*signed(FMAP_70_38);
			MULT_39(69)<=signed(DIN_39_7)*signed(FMAP_70_39);
			MULT_40(69)<=signed(DIN_40_7)*signed(FMAP_70_40);
			MULT_41(69)<=signed(DIN_41_7)*signed(FMAP_70_41);
			MULT_42(69)<=signed(DIN_42_7)*signed(FMAP_70_42);
			MULT_43(69)<=signed(DIN_43_7)*signed(FMAP_70_43);
			MULT_44(69)<=signed(DIN_44_7)*signed(FMAP_70_44);
			MULT_45(69)<=signed(DIN_45_7)*signed(FMAP_70_45);
			MULT_46(69)<=signed(DIN_46_7)*signed(FMAP_70_46);
			MULT_47(69)<=signed(DIN_47_7)*signed(FMAP_70_47);
			MULT_48(69)<=signed(DIN_48_7)*signed(FMAP_70_48);
			MULT_49(69)<=signed(DIN_49_7)*signed(FMAP_70_49);
			MULT_50(69)<=signed(DIN_50_7)*signed(FMAP_70_50);
			MULT_51(69)<=signed(DIN_51_7)*signed(FMAP_70_51);
			MULT_52(69)<=signed(DIN_52_7)*signed(FMAP_70_52);
			MULT_53(69)<=signed(DIN_53_7)*signed(FMAP_70_53);
			MULT_54(69)<=signed(DIN_54_7)*signed(FMAP_70_54);
			MULT_55(69)<=signed(DIN_55_7)*signed(FMAP_70_55);
			MULT_56(69)<=signed(DIN_56_7)*signed(FMAP_70_56);
			MULT_57(69)<=signed(DIN_57_7)*signed(FMAP_70_57);
			MULT_58(69)<=signed(DIN_58_7)*signed(FMAP_70_58);
			MULT_59(69)<=signed(DIN_59_7)*signed(FMAP_70_59);
			MULT_60(69)<=signed(DIN_60_7)*signed(FMAP_70_60);
			MULT_61(69)<=signed(DIN_61_7)*signed(FMAP_70_61);
			MULT_62(69)<=signed(DIN_62_7)*signed(FMAP_70_62);
			MULT_63(69)<=signed(DIN_63_7)*signed(FMAP_70_63);
			MULT_64(69)<=signed(DIN_64_7)*signed(FMAP_70_64);
			MULT_65(69)<=signed(DIN_65_7)*signed(FMAP_70_65);
			MULT_66(69)<=signed(DIN_66_7)*signed(FMAP_70_66);
			MULT_67(69)<=signed(DIN_67_7)*signed(FMAP_70_67);
			MULT_68(69)<=signed(DIN_68_7)*signed(FMAP_70_68);
			MULT_69(69)<=signed(DIN_69_7)*signed(FMAP_70_69);
			MULT_70(69)<=signed(DIN_70_7)*signed(FMAP_70_70);
			MULT_71(69)<=signed(DIN_71_7)*signed(FMAP_70_71);
			MULT_72(69)<=signed(DIN_72_7)*signed(FMAP_70_72);
			MULT_73(69)<=signed(DIN_73_7)*signed(FMAP_70_73);
			MULT_74(69)<=signed(DIN_74_7)*signed(FMAP_70_74);
			MULT_75(69)<=signed(DIN_75_7)*signed(FMAP_70_75);
			MULT_76(69)<=signed(DIN_76_7)*signed(FMAP_70_76);
			MULT_77(69)<=signed(DIN_77_7)*signed(FMAP_70_77);
			MULT_78(69)<=signed(DIN_78_7)*signed(FMAP_70_78);
			MULT_79(69)<=signed(DIN_79_7)*signed(FMAP_70_79);
			MULT_80(69)<=signed(DIN_80_7)*signed(FMAP_70_80);
			MULT_81(69)<=signed(DIN_81_7)*signed(FMAP_70_81);
			MULT_82(69)<=signed(DIN_82_7)*signed(FMAP_70_82);
			MULT_83(69)<=signed(DIN_83_7)*signed(FMAP_70_83);
			MULT_84(69)<=signed(DIN_84_7)*signed(FMAP_70_84);
			MULT_85(69)<=signed(DIN_85_7)*signed(FMAP_70_85);
			MULT_86(69)<=signed(DIN_86_7)*signed(FMAP_70_86);
			MULT_87(69)<=signed(DIN_87_7)*signed(FMAP_70_87);
			MULT_88(69)<=signed(DIN_88_7)*signed(FMAP_70_88);
			MULT_89(69)<=signed(DIN_89_7)*signed(FMAP_70_89);
			MULT_90(69)<=signed(DIN_90_7)*signed(FMAP_70_90);
			MULT_91(69)<=signed(DIN_91_7)*signed(FMAP_70_91);
			MULT_92(69)<=signed(DIN_92_7)*signed(FMAP_70_92);
			MULT_93(69)<=signed(DIN_93_7)*signed(FMAP_70_93);
			MULT_94(69)<=signed(DIN_94_7)*signed(FMAP_70_94);
			MULT_95(69)<=signed(DIN_95_7)*signed(FMAP_70_95);
			MULT_96(69)<=signed(DIN_96_7)*signed(FMAP_70_96);
			MULT_97(69)<=signed(DIN_97_7)*signed(FMAP_70_97);
			MULT_98(69)<=signed(DIN_98_7)*signed(FMAP_70_98);
			MULT_99(69)<=signed(DIN_99_7)*signed(FMAP_70_99);
			MULT_100(69)<=signed(DIN_100_7)*signed(FMAP_70_100);
			MULT_101(69)<=signed(DIN_101_7)*signed(FMAP_70_101);
			MULT_102(69)<=signed(DIN_102_7)*signed(FMAP_70_102);
			MULT_103(69)<=signed(DIN_103_7)*signed(FMAP_70_103);
			MULT_104(69)<=signed(DIN_104_7)*signed(FMAP_70_104);
			MULT_105(69)<=signed(DIN_105_7)*signed(FMAP_70_105);
			MULT_106(69)<=signed(DIN_106_7)*signed(FMAP_70_106);
			MULT_107(69)<=signed(DIN_107_7)*signed(FMAP_70_107);
			MULT_108(69)<=signed(DIN_108_7)*signed(FMAP_70_108);
			MULT_109(69)<=signed(DIN_109_7)*signed(FMAP_70_109);
			MULT_110(69)<=signed(DIN_110_7)*signed(FMAP_70_110);
			MULT_111(69)<=signed(DIN_111_7)*signed(FMAP_70_111);
			MULT_112(69)<=signed(DIN_112_7)*signed(FMAP_70_112);
			MULT_113(69)<=signed(DIN_113_7)*signed(FMAP_70_113);
			MULT_114(69)<=signed(DIN_114_7)*signed(FMAP_70_114);
			MULT_115(69)<=signed(DIN_115_7)*signed(FMAP_70_115);
			MULT_116(69)<=signed(DIN_116_7)*signed(FMAP_70_116);
			MULT_117(69)<=signed(DIN_117_7)*signed(FMAP_70_117);
			MULT_118(69)<=signed(DIN_118_7)*signed(FMAP_70_118);
			MULT_119(69)<=signed(DIN_119_7)*signed(FMAP_70_119);
			MULT_120(69)<=signed(DIN_120_7)*signed(FMAP_70_120);

			MULT_1(70)<=signed(DIN_1_7)*signed(FMAP_71_1);
			MULT_2(70)<=signed(DIN_2_7)*signed(FMAP_71_2);
			MULT_3(70)<=signed(DIN_3_7)*signed(FMAP_71_3);
			MULT_4(70)<=signed(DIN_4_7)*signed(FMAP_71_4);
			MULT_5(70)<=signed(DIN_5_7)*signed(FMAP_71_5);
			MULT_6(70)<=signed(DIN_6_7)*signed(FMAP_71_6);
			MULT_7(70)<=signed(DIN_7_7)*signed(FMAP_71_7);
			MULT_8(70)<=signed(DIN_8_7)*signed(FMAP_71_8);
			MULT_9(70)<=signed(DIN_9_7)*signed(FMAP_71_9);
			MULT_10(70)<=signed(DIN_10_7)*signed(FMAP_71_10);
			MULT_11(70)<=signed(DIN_11_7)*signed(FMAP_71_11);
			MULT_12(70)<=signed(DIN_12_7)*signed(FMAP_71_12);
			MULT_13(70)<=signed(DIN_13_7)*signed(FMAP_71_13);
			MULT_14(70)<=signed(DIN_14_7)*signed(FMAP_71_14);
			MULT_15(70)<=signed(DIN_15_7)*signed(FMAP_71_15);
			MULT_16(70)<=signed(DIN_16_7)*signed(FMAP_71_16);
			MULT_17(70)<=signed(DIN_17_7)*signed(FMAP_71_17);
			MULT_18(70)<=signed(DIN_18_7)*signed(FMAP_71_18);
			MULT_19(70)<=signed(DIN_19_7)*signed(FMAP_71_19);
			MULT_20(70)<=signed(DIN_20_7)*signed(FMAP_71_20);
			MULT_21(70)<=signed(DIN_21_7)*signed(FMAP_71_21);
			MULT_22(70)<=signed(DIN_22_7)*signed(FMAP_71_22);
			MULT_23(70)<=signed(DIN_23_7)*signed(FMAP_71_23);
			MULT_24(70)<=signed(DIN_24_7)*signed(FMAP_71_24);
			MULT_25(70)<=signed(DIN_25_7)*signed(FMAP_71_25);
			MULT_26(70)<=signed(DIN_26_7)*signed(FMAP_71_26);
			MULT_27(70)<=signed(DIN_27_7)*signed(FMAP_71_27);
			MULT_28(70)<=signed(DIN_28_7)*signed(FMAP_71_28);
			MULT_29(70)<=signed(DIN_29_7)*signed(FMAP_71_29);
			MULT_30(70)<=signed(DIN_30_7)*signed(FMAP_71_30);
			MULT_31(70)<=signed(DIN_31_7)*signed(FMAP_71_31);
			MULT_32(70)<=signed(DIN_32_7)*signed(FMAP_71_32);
			MULT_33(70)<=signed(DIN_33_7)*signed(FMAP_71_33);
			MULT_34(70)<=signed(DIN_34_7)*signed(FMAP_71_34);
			MULT_35(70)<=signed(DIN_35_7)*signed(FMAP_71_35);
			MULT_36(70)<=signed(DIN_36_7)*signed(FMAP_71_36);
			MULT_37(70)<=signed(DIN_37_7)*signed(FMAP_71_37);
			MULT_38(70)<=signed(DIN_38_7)*signed(FMAP_71_38);
			MULT_39(70)<=signed(DIN_39_7)*signed(FMAP_71_39);
			MULT_40(70)<=signed(DIN_40_7)*signed(FMAP_71_40);
			MULT_41(70)<=signed(DIN_41_7)*signed(FMAP_71_41);
			MULT_42(70)<=signed(DIN_42_7)*signed(FMAP_71_42);
			MULT_43(70)<=signed(DIN_43_7)*signed(FMAP_71_43);
			MULT_44(70)<=signed(DIN_44_7)*signed(FMAP_71_44);
			MULT_45(70)<=signed(DIN_45_7)*signed(FMAP_71_45);
			MULT_46(70)<=signed(DIN_46_7)*signed(FMAP_71_46);
			MULT_47(70)<=signed(DIN_47_7)*signed(FMAP_71_47);
			MULT_48(70)<=signed(DIN_48_7)*signed(FMAP_71_48);
			MULT_49(70)<=signed(DIN_49_7)*signed(FMAP_71_49);
			MULT_50(70)<=signed(DIN_50_7)*signed(FMAP_71_50);
			MULT_51(70)<=signed(DIN_51_7)*signed(FMAP_71_51);
			MULT_52(70)<=signed(DIN_52_7)*signed(FMAP_71_52);
			MULT_53(70)<=signed(DIN_53_7)*signed(FMAP_71_53);
			MULT_54(70)<=signed(DIN_54_7)*signed(FMAP_71_54);
			MULT_55(70)<=signed(DIN_55_7)*signed(FMAP_71_55);
			MULT_56(70)<=signed(DIN_56_7)*signed(FMAP_71_56);
			MULT_57(70)<=signed(DIN_57_7)*signed(FMAP_71_57);
			MULT_58(70)<=signed(DIN_58_7)*signed(FMAP_71_58);
			MULT_59(70)<=signed(DIN_59_7)*signed(FMAP_71_59);
			MULT_60(70)<=signed(DIN_60_7)*signed(FMAP_71_60);
			MULT_61(70)<=signed(DIN_61_7)*signed(FMAP_71_61);
			MULT_62(70)<=signed(DIN_62_7)*signed(FMAP_71_62);
			MULT_63(70)<=signed(DIN_63_7)*signed(FMAP_71_63);
			MULT_64(70)<=signed(DIN_64_7)*signed(FMAP_71_64);
			MULT_65(70)<=signed(DIN_65_7)*signed(FMAP_71_65);
			MULT_66(70)<=signed(DIN_66_7)*signed(FMAP_71_66);
			MULT_67(70)<=signed(DIN_67_7)*signed(FMAP_71_67);
			MULT_68(70)<=signed(DIN_68_7)*signed(FMAP_71_68);
			MULT_69(70)<=signed(DIN_69_7)*signed(FMAP_71_69);
			MULT_70(70)<=signed(DIN_70_7)*signed(FMAP_71_70);
			MULT_71(70)<=signed(DIN_71_7)*signed(FMAP_71_71);
			MULT_72(70)<=signed(DIN_72_7)*signed(FMAP_71_72);
			MULT_73(70)<=signed(DIN_73_7)*signed(FMAP_71_73);
			MULT_74(70)<=signed(DIN_74_7)*signed(FMAP_71_74);
			MULT_75(70)<=signed(DIN_75_7)*signed(FMAP_71_75);
			MULT_76(70)<=signed(DIN_76_7)*signed(FMAP_71_76);
			MULT_77(70)<=signed(DIN_77_7)*signed(FMAP_71_77);
			MULT_78(70)<=signed(DIN_78_7)*signed(FMAP_71_78);
			MULT_79(70)<=signed(DIN_79_7)*signed(FMAP_71_79);
			MULT_80(70)<=signed(DIN_80_7)*signed(FMAP_71_80);
			MULT_81(70)<=signed(DIN_81_7)*signed(FMAP_71_81);
			MULT_82(70)<=signed(DIN_82_7)*signed(FMAP_71_82);
			MULT_83(70)<=signed(DIN_83_7)*signed(FMAP_71_83);
			MULT_84(70)<=signed(DIN_84_7)*signed(FMAP_71_84);
			MULT_85(70)<=signed(DIN_85_7)*signed(FMAP_71_85);
			MULT_86(70)<=signed(DIN_86_7)*signed(FMAP_71_86);
			MULT_87(70)<=signed(DIN_87_7)*signed(FMAP_71_87);
			MULT_88(70)<=signed(DIN_88_7)*signed(FMAP_71_88);
			MULT_89(70)<=signed(DIN_89_7)*signed(FMAP_71_89);
			MULT_90(70)<=signed(DIN_90_7)*signed(FMAP_71_90);
			MULT_91(70)<=signed(DIN_91_7)*signed(FMAP_71_91);
			MULT_92(70)<=signed(DIN_92_7)*signed(FMAP_71_92);
			MULT_93(70)<=signed(DIN_93_7)*signed(FMAP_71_93);
			MULT_94(70)<=signed(DIN_94_7)*signed(FMAP_71_94);
			MULT_95(70)<=signed(DIN_95_7)*signed(FMAP_71_95);
			MULT_96(70)<=signed(DIN_96_7)*signed(FMAP_71_96);
			MULT_97(70)<=signed(DIN_97_7)*signed(FMAP_71_97);
			MULT_98(70)<=signed(DIN_98_7)*signed(FMAP_71_98);
			MULT_99(70)<=signed(DIN_99_7)*signed(FMAP_71_99);
			MULT_100(70)<=signed(DIN_100_7)*signed(FMAP_71_100);
			MULT_101(70)<=signed(DIN_101_7)*signed(FMAP_71_101);
			MULT_102(70)<=signed(DIN_102_7)*signed(FMAP_71_102);
			MULT_103(70)<=signed(DIN_103_7)*signed(FMAP_71_103);
			MULT_104(70)<=signed(DIN_104_7)*signed(FMAP_71_104);
			MULT_105(70)<=signed(DIN_105_7)*signed(FMAP_71_105);
			MULT_106(70)<=signed(DIN_106_7)*signed(FMAP_71_106);
			MULT_107(70)<=signed(DIN_107_7)*signed(FMAP_71_107);
			MULT_108(70)<=signed(DIN_108_7)*signed(FMAP_71_108);
			MULT_109(70)<=signed(DIN_109_7)*signed(FMAP_71_109);
			MULT_110(70)<=signed(DIN_110_7)*signed(FMAP_71_110);
			MULT_111(70)<=signed(DIN_111_7)*signed(FMAP_71_111);
			MULT_112(70)<=signed(DIN_112_7)*signed(FMAP_71_112);
			MULT_113(70)<=signed(DIN_113_7)*signed(FMAP_71_113);
			MULT_114(70)<=signed(DIN_114_7)*signed(FMAP_71_114);
			MULT_115(70)<=signed(DIN_115_7)*signed(FMAP_71_115);
			MULT_116(70)<=signed(DIN_116_7)*signed(FMAP_71_116);
			MULT_117(70)<=signed(DIN_117_7)*signed(FMAP_71_117);
			MULT_118(70)<=signed(DIN_118_7)*signed(FMAP_71_118);
			MULT_119(70)<=signed(DIN_119_7)*signed(FMAP_71_119);
			MULT_120(70)<=signed(DIN_120_7)*signed(FMAP_71_120);

			MULT_1(71)<=signed(DIN_1_7)*signed(FMAP_72_1);
			MULT_2(71)<=signed(DIN_2_7)*signed(FMAP_72_2);
			MULT_3(71)<=signed(DIN_3_7)*signed(FMAP_72_3);
			MULT_4(71)<=signed(DIN_4_7)*signed(FMAP_72_4);
			MULT_5(71)<=signed(DIN_5_7)*signed(FMAP_72_5);
			MULT_6(71)<=signed(DIN_6_7)*signed(FMAP_72_6);
			MULT_7(71)<=signed(DIN_7_7)*signed(FMAP_72_7);
			MULT_8(71)<=signed(DIN_8_7)*signed(FMAP_72_8);
			MULT_9(71)<=signed(DIN_9_7)*signed(FMAP_72_9);
			MULT_10(71)<=signed(DIN_10_7)*signed(FMAP_72_10);
			MULT_11(71)<=signed(DIN_11_7)*signed(FMAP_72_11);
			MULT_12(71)<=signed(DIN_12_7)*signed(FMAP_72_12);
			MULT_13(71)<=signed(DIN_13_7)*signed(FMAP_72_13);
			MULT_14(71)<=signed(DIN_14_7)*signed(FMAP_72_14);
			MULT_15(71)<=signed(DIN_15_7)*signed(FMAP_72_15);
			MULT_16(71)<=signed(DIN_16_7)*signed(FMAP_72_16);
			MULT_17(71)<=signed(DIN_17_7)*signed(FMAP_72_17);
			MULT_18(71)<=signed(DIN_18_7)*signed(FMAP_72_18);
			MULT_19(71)<=signed(DIN_19_7)*signed(FMAP_72_19);
			MULT_20(71)<=signed(DIN_20_7)*signed(FMAP_72_20);
			MULT_21(71)<=signed(DIN_21_7)*signed(FMAP_72_21);
			MULT_22(71)<=signed(DIN_22_7)*signed(FMAP_72_22);
			MULT_23(71)<=signed(DIN_23_7)*signed(FMAP_72_23);
			MULT_24(71)<=signed(DIN_24_7)*signed(FMAP_72_24);
			MULT_25(71)<=signed(DIN_25_7)*signed(FMAP_72_25);
			MULT_26(71)<=signed(DIN_26_7)*signed(FMAP_72_26);
			MULT_27(71)<=signed(DIN_27_7)*signed(FMAP_72_27);
			MULT_28(71)<=signed(DIN_28_7)*signed(FMAP_72_28);
			MULT_29(71)<=signed(DIN_29_7)*signed(FMAP_72_29);
			MULT_30(71)<=signed(DIN_30_7)*signed(FMAP_72_30);
			MULT_31(71)<=signed(DIN_31_7)*signed(FMAP_72_31);
			MULT_32(71)<=signed(DIN_32_7)*signed(FMAP_72_32);
			MULT_33(71)<=signed(DIN_33_7)*signed(FMAP_72_33);
			MULT_34(71)<=signed(DIN_34_7)*signed(FMAP_72_34);
			MULT_35(71)<=signed(DIN_35_7)*signed(FMAP_72_35);
			MULT_36(71)<=signed(DIN_36_7)*signed(FMAP_72_36);
			MULT_37(71)<=signed(DIN_37_7)*signed(FMAP_72_37);
			MULT_38(71)<=signed(DIN_38_7)*signed(FMAP_72_38);
			MULT_39(71)<=signed(DIN_39_7)*signed(FMAP_72_39);
			MULT_40(71)<=signed(DIN_40_7)*signed(FMAP_72_40);
			MULT_41(71)<=signed(DIN_41_7)*signed(FMAP_72_41);
			MULT_42(71)<=signed(DIN_42_7)*signed(FMAP_72_42);
			MULT_43(71)<=signed(DIN_43_7)*signed(FMAP_72_43);
			MULT_44(71)<=signed(DIN_44_7)*signed(FMAP_72_44);
			MULT_45(71)<=signed(DIN_45_7)*signed(FMAP_72_45);
			MULT_46(71)<=signed(DIN_46_7)*signed(FMAP_72_46);
			MULT_47(71)<=signed(DIN_47_7)*signed(FMAP_72_47);
			MULT_48(71)<=signed(DIN_48_7)*signed(FMAP_72_48);
			MULT_49(71)<=signed(DIN_49_7)*signed(FMAP_72_49);
			MULT_50(71)<=signed(DIN_50_7)*signed(FMAP_72_50);
			MULT_51(71)<=signed(DIN_51_7)*signed(FMAP_72_51);
			MULT_52(71)<=signed(DIN_52_7)*signed(FMAP_72_52);
			MULT_53(71)<=signed(DIN_53_7)*signed(FMAP_72_53);
			MULT_54(71)<=signed(DIN_54_7)*signed(FMAP_72_54);
			MULT_55(71)<=signed(DIN_55_7)*signed(FMAP_72_55);
			MULT_56(71)<=signed(DIN_56_7)*signed(FMAP_72_56);
			MULT_57(71)<=signed(DIN_57_7)*signed(FMAP_72_57);
			MULT_58(71)<=signed(DIN_58_7)*signed(FMAP_72_58);
			MULT_59(71)<=signed(DIN_59_7)*signed(FMAP_72_59);
			MULT_60(71)<=signed(DIN_60_7)*signed(FMAP_72_60);
			MULT_61(71)<=signed(DIN_61_7)*signed(FMAP_72_61);
			MULT_62(71)<=signed(DIN_62_7)*signed(FMAP_72_62);
			MULT_63(71)<=signed(DIN_63_7)*signed(FMAP_72_63);
			MULT_64(71)<=signed(DIN_64_7)*signed(FMAP_72_64);
			MULT_65(71)<=signed(DIN_65_7)*signed(FMAP_72_65);
			MULT_66(71)<=signed(DIN_66_7)*signed(FMAP_72_66);
			MULT_67(71)<=signed(DIN_67_7)*signed(FMAP_72_67);
			MULT_68(71)<=signed(DIN_68_7)*signed(FMAP_72_68);
			MULT_69(71)<=signed(DIN_69_7)*signed(FMAP_72_69);
			MULT_70(71)<=signed(DIN_70_7)*signed(FMAP_72_70);
			MULT_71(71)<=signed(DIN_71_7)*signed(FMAP_72_71);
			MULT_72(71)<=signed(DIN_72_7)*signed(FMAP_72_72);
			MULT_73(71)<=signed(DIN_73_7)*signed(FMAP_72_73);
			MULT_74(71)<=signed(DIN_74_7)*signed(FMAP_72_74);
			MULT_75(71)<=signed(DIN_75_7)*signed(FMAP_72_75);
			MULT_76(71)<=signed(DIN_76_7)*signed(FMAP_72_76);
			MULT_77(71)<=signed(DIN_77_7)*signed(FMAP_72_77);
			MULT_78(71)<=signed(DIN_78_7)*signed(FMAP_72_78);
			MULT_79(71)<=signed(DIN_79_7)*signed(FMAP_72_79);
			MULT_80(71)<=signed(DIN_80_7)*signed(FMAP_72_80);
			MULT_81(71)<=signed(DIN_81_7)*signed(FMAP_72_81);
			MULT_82(71)<=signed(DIN_82_7)*signed(FMAP_72_82);
			MULT_83(71)<=signed(DIN_83_7)*signed(FMAP_72_83);
			MULT_84(71)<=signed(DIN_84_7)*signed(FMAP_72_84);
			MULT_85(71)<=signed(DIN_85_7)*signed(FMAP_72_85);
			MULT_86(71)<=signed(DIN_86_7)*signed(FMAP_72_86);
			MULT_87(71)<=signed(DIN_87_7)*signed(FMAP_72_87);
			MULT_88(71)<=signed(DIN_88_7)*signed(FMAP_72_88);
			MULT_89(71)<=signed(DIN_89_7)*signed(FMAP_72_89);
			MULT_90(71)<=signed(DIN_90_7)*signed(FMAP_72_90);
			MULT_91(71)<=signed(DIN_91_7)*signed(FMAP_72_91);
			MULT_92(71)<=signed(DIN_92_7)*signed(FMAP_72_92);
			MULT_93(71)<=signed(DIN_93_7)*signed(FMAP_72_93);
			MULT_94(71)<=signed(DIN_94_7)*signed(FMAP_72_94);
			MULT_95(71)<=signed(DIN_95_7)*signed(FMAP_72_95);
			MULT_96(71)<=signed(DIN_96_7)*signed(FMAP_72_96);
			MULT_97(71)<=signed(DIN_97_7)*signed(FMAP_72_97);
			MULT_98(71)<=signed(DIN_98_7)*signed(FMAP_72_98);
			MULT_99(71)<=signed(DIN_99_7)*signed(FMAP_72_99);
			MULT_100(71)<=signed(DIN_100_7)*signed(FMAP_72_100);
			MULT_101(71)<=signed(DIN_101_7)*signed(FMAP_72_101);
			MULT_102(71)<=signed(DIN_102_7)*signed(FMAP_72_102);
			MULT_103(71)<=signed(DIN_103_7)*signed(FMAP_72_103);
			MULT_104(71)<=signed(DIN_104_7)*signed(FMAP_72_104);
			MULT_105(71)<=signed(DIN_105_7)*signed(FMAP_72_105);
			MULT_106(71)<=signed(DIN_106_7)*signed(FMAP_72_106);
			MULT_107(71)<=signed(DIN_107_7)*signed(FMAP_72_107);
			MULT_108(71)<=signed(DIN_108_7)*signed(FMAP_72_108);
			MULT_109(71)<=signed(DIN_109_7)*signed(FMAP_72_109);
			MULT_110(71)<=signed(DIN_110_7)*signed(FMAP_72_110);
			MULT_111(71)<=signed(DIN_111_7)*signed(FMAP_72_111);
			MULT_112(71)<=signed(DIN_112_7)*signed(FMAP_72_112);
			MULT_113(71)<=signed(DIN_113_7)*signed(FMAP_72_113);
			MULT_114(71)<=signed(DIN_114_7)*signed(FMAP_72_114);
			MULT_115(71)<=signed(DIN_115_7)*signed(FMAP_72_115);
			MULT_116(71)<=signed(DIN_116_7)*signed(FMAP_72_116);
			MULT_117(71)<=signed(DIN_117_7)*signed(FMAP_72_117);
			MULT_118(71)<=signed(DIN_118_7)*signed(FMAP_72_118);
			MULT_119(71)<=signed(DIN_119_7)*signed(FMAP_72_119);
			MULT_120(71)<=signed(DIN_120_7)*signed(FMAP_72_120);

			MULT_1(72)<=signed(DIN_1_7)*signed(FMAP_73_1);
			MULT_2(72)<=signed(DIN_2_7)*signed(FMAP_73_2);
			MULT_3(72)<=signed(DIN_3_7)*signed(FMAP_73_3);
			MULT_4(72)<=signed(DIN_4_7)*signed(FMAP_73_4);
			MULT_5(72)<=signed(DIN_5_7)*signed(FMAP_73_5);
			MULT_6(72)<=signed(DIN_6_7)*signed(FMAP_73_6);
			MULT_7(72)<=signed(DIN_7_7)*signed(FMAP_73_7);
			MULT_8(72)<=signed(DIN_8_7)*signed(FMAP_73_8);
			MULT_9(72)<=signed(DIN_9_7)*signed(FMAP_73_9);
			MULT_10(72)<=signed(DIN_10_7)*signed(FMAP_73_10);
			MULT_11(72)<=signed(DIN_11_7)*signed(FMAP_73_11);
			MULT_12(72)<=signed(DIN_12_7)*signed(FMAP_73_12);
			MULT_13(72)<=signed(DIN_13_7)*signed(FMAP_73_13);
			MULT_14(72)<=signed(DIN_14_7)*signed(FMAP_73_14);
			MULT_15(72)<=signed(DIN_15_7)*signed(FMAP_73_15);
			MULT_16(72)<=signed(DIN_16_7)*signed(FMAP_73_16);
			MULT_17(72)<=signed(DIN_17_7)*signed(FMAP_73_17);
			MULT_18(72)<=signed(DIN_18_7)*signed(FMAP_73_18);
			MULT_19(72)<=signed(DIN_19_7)*signed(FMAP_73_19);
			MULT_20(72)<=signed(DIN_20_7)*signed(FMAP_73_20);
			MULT_21(72)<=signed(DIN_21_7)*signed(FMAP_73_21);
			MULT_22(72)<=signed(DIN_22_7)*signed(FMAP_73_22);
			MULT_23(72)<=signed(DIN_23_7)*signed(FMAP_73_23);
			MULT_24(72)<=signed(DIN_24_7)*signed(FMAP_73_24);
			MULT_25(72)<=signed(DIN_25_7)*signed(FMAP_73_25);
			MULT_26(72)<=signed(DIN_26_7)*signed(FMAP_73_26);
			MULT_27(72)<=signed(DIN_27_7)*signed(FMAP_73_27);
			MULT_28(72)<=signed(DIN_28_7)*signed(FMAP_73_28);
			MULT_29(72)<=signed(DIN_29_7)*signed(FMAP_73_29);
			MULT_30(72)<=signed(DIN_30_7)*signed(FMAP_73_30);
			MULT_31(72)<=signed(DIN_31_7)*signed(FMAP_73_31);
			MULT_32(72)<=signed(DIN_32_7)*signed(FMAP_73_32);
			MULT_33(72)<=signed(DIN_33_7)*signed(FMAP_73_33);
			MULT_34(72)<=signed(DIN_34_7)*signed(FMAP_73_34);
			MULT_35(72)<=signed(DIN_35_7)*signed(FMAP_73_35);
			MULT_36(72)<=signed(DIN_36_7)*signed(FMAP_73_36);
			MULT_37(72)<=signed(DIN_37_7)*signed(FMAP_73_37);
			MULT_38(72)<=signed(DIN_38_7)*signed(FMAP_73_38);
			MULT_39(72)<=signed(DIN_39_7)*signed(FMAP_73_39);
			MULT_40(72)<=signed(DIN_40_7)*signed(FMAP_73_40);
			MULT_41(72)<=signed(DIN_41_7)*signed(FMAP_73_41);
			MULT_42(72)<=signed(DIN_42_7)*signed(FMAP_73_42);
			MULT_43(72)<=signed(DIN_43_7)*signed(FMAP_73_43);
			MULT_44(72)<=signed(DIN_44_7)*signed(FMAP_73_44);
			MULT_45(72)<=signed(DIN_45_7)*signed(FMAP_73_45);
			MULT_46(72)<=signed(DIN_46_7)*signed(FMAP_73_46);
			MULT_47(72)<=signed(DIN_47_7)*signed(FMAP_73_47);
			MULT_48(72)<=signed(DIN_48_7)*signed(FMAP_73_48);
			MULT_49(72)<=signed(DIN_49_7)*signed(FMAP_73_49);
			MULT_50(72)<=signed(DIN_50_7)*signed(FMAP_73_50);
			MULT_51(72)<=signed(DIN_51_7)*signed(FMAP_73_51);
			MULT_52(72)<=signed(DIN_52_7)*signed(FMAP_73_52);
			MULT_53(72)<=signed(DIN_53_7)*signed(FMAP_73_53);
			MULT_54(72)<=signed(DIN_54_7)*signed(FMAP_73_54);
			MULT_55(72)<=signed(DIN_55_7)*signed(FMAP_73_55);
			MULT_56(72)<=signed(DIN_56_7)*signed(FMAP_73_56);
			MULT_57(72)<=signed(DIN_57_7)*signed(FMAP_73_57);
			MULT_58(72)<=signed(DIN_58_7)*signed(FMAP_73_58);
			MULT_59(72)<=signed(DIN_59_7)*signed(FMAP_73_59);
			MULT_60(72)<=signed(DIN_60_7)*signed(FMAP_73_60);
			MULT_61(72)<=signed(DIN_61_7)*signed(FMAP_73_61);
			MULT_62(72)<=signed(DIN_62_7)*signed(FMAP_73_62);
			MULT_63(72)<=signed(DIN_63_7)*signed(FMAP_73_63);
			MULT_64(72)<=signed(DIN_64_7)*signed(FMAP_73_64);
			MULT_65(72)<=signed(DIN_65_7)*signed(FMAP_73_65);
			MULT_66(72)<=signed(DIN_66_7)*signed(FMAP_73_66);
			MULT_67(72)<=signed(DIN_67_7)*signed(FMAP_73_67);
			MULT_68(72)<=signed(DIN_68_7)*signed(FMAP_73_68);
			MULT_69(72)<=signed(DIN_69_7)*signed(FMAP_73_69);
			MULT_70(72)<=signed(DIN_70_7)*signed(FMAP_73_70);
			MULT_71(72)<=signed(DIN_71_7)*signed(FMAP_73_71);
			MULT_72(72)<=signed(DIN_72_7)*signed(FMAP_73_72);
			MULT_73(72)<=signed(DIN_73_7)*signed(FMAP_73_73);
			MULT_74(72)<=signed(DIN_74_7)*signed(FMAP_73_74);
			MULT_75(72)<=signed(DIN_75_7)*signed(FMAP_73_75);
			MULT_76(72)<=signed(DIN_76_7)*signed(FMAP_73_76);
			MULT_77(72)<=signed(DIN_77_7)*signed(FMAP_73_77);
			MULT_78(72)<=signed(DIN_78_7)*signed(FMAP_73_78);
			MULT_79(72)<=signed(DIN_79_7)*signed(FMAP_73_79);
			MULT_80(72)<=signed(DIN_80_7)*signed(FMAP_73_80);
			MULT_81(72)<=signed(DIN_81_7)*signed(FMAP_73_81);
			MULT_82(72)<=signed(DIN_82_7)*signed(FMAP_73_82);
			MULT_83(72)<=signed(DIN_83_7)*signed(FMAP_73_83);
			MULT_84(72)<=signed(DIN_84_7)*signed(FMAP_73_84);
			MULT_85(72)<=signed(DIN_85_7)*signed(FMAP_73_85);
			MULT_86(72)<=signed(DIN_86_7)*signed(FMAP_73_86);
			MULT_87(72)<=signed(DIN_87_7)*signed(FMAP_73_87);
			MULT_88(72)<=signed(DIN_88_7)*signed(FMAP_73_88);
			MULT_89(72)<=signed(DIN_89_7)*signed(FMAP_73_89);
			MULT_90(72)<=signed(DIN_90_7)*signed(FMAP_73_90);
			MULT_91(72)<=signed(DIN_91_7)*signed(FMAP_73_91);
			MULT_92(72)<=signed(DIN_92_7)*signed(FMAP_73_92);
			MULT_93(72)<=signed(DIN_93_7)*signed(FMAP_73_93);
			MULT_94(72)<=signed(DIN_94_7)*signed(FMAP_73_94);
			MULT_95(72)<=signed(DIN_95_7)*signed(FMAP_73_95);
			MULT_96(72)<=signed(DIN_96_7)*signed(FMAP_73_96);
			MULT_97(72)<=signed(DIN_97_7)*signed(FMAP_73_97);
			MULT_98(72)<=signed(DIN_98_7)*signed(FMAP_73_98);
			MULT_99(72)<=signed(DIN_99_7)*signed(FMAP_73_99);
			MULT_100(72)<=signed(DIN_100_7)*signed(FMAP_73_100);
			MULT_101(72)<=signed(DIN_101_7)*signed(FMAP_73_101);
			MULT_102(72)<=signed(DIN_102_7)*signed(FMAP_73_102);
			MULT_103(72)<=signed(DIN_103_7)*signed(FMAP_73_103);
			MULT_104(72)<=signed(DIN_104_7)*signed(FMAP_73_104);
			MULT_105(72)<=signed(DIN_105_7)*signed(FMAP_73_105);
			MULT_106(72)<=signed(DIN_106_7)*signed(FMAP_73_106);
			MULT_107(72)<=signed(DIN_107_7)*signed(FMAP_73_107);
			MULT_108(72)<=signed(DIN_108_7)*signed(FMAP_73_108);
			MULT_109(72)<=signed(DIN_109_7)*signed(FMAP_73_109);
			MULT_110(72)<=signed(DIN_110_7)*signed(FMAP_73_110);
			MULT_111(72)<=signed(DIN_111_7)*signed(FMAP_73_111);
			MULT_112(72)<=signed(DIN_112_7)*signed(FMAP_73_112);
			MULT_113(72)<=signed(DIN_113_7)*signed(FMAP_73_113);
			MULT_114(72)<=signed(DIN_114_7)*signed(FMAP_73_114);
			MULT_115(72)<=signed(DIN_115_7)*signed(FMAP_73_115);
			MULT_116(72)<=signed(DIN_116_7)*signed(FMAP_73_116);
			MULT_117(72)<=signed(DIN_117_7)*signed(FMAP_73_117);
			MULT_118(72)<=signed(DIN_118_7)*signed(FMAP_73_118);
			MULT_119(72)<=signed(DIN_119_7)*signed(FMAP_73_119);
			MULT_120(72)<=signed(DIN_120_7)*signed(FMAP_73_120);

			MULT_1(73)<=signed(DIN_1_7)*signed(FMAP_74_1);
			MULT_2(73)<=signed(DIN_2_7)*signed(FMAP_74_2);
			MULT_3(73)<=signed(DIN_3_7)*signed(FMAP_74_3);
			MULT_4(73)<=signed(DIN_4_7)*signed(FMAP_74_4);
			MULT_5(73)<=signed(DIN_5_7)*signed(FMAP_74_5);
			MULT_6(73)<=signed(DIN_6_7)*signed(FMAP_74_6);
			MULT_7(73)<=signed(DIN_7_7)*signed(FMAP_74_7);
			MULT_8(73)<=signed(DIN_8_7)*signed(FMAP_74_8);
			MULT_9(73)<=signed(DIN_9_7)*signed(FMAP_74_9);
			MULT_10(73)<=signed(DIN_10_7)*signed(FMAP_74_10);
			MULT_11(73)<=signed(DIN_11_7)*signed(FMAP_74_11);
			MULT_12(73)<=signed(DIN_12_7)*signed(FMAP_74_12);
			MULT_13(73)<=signed(DIN_13_7)*signed(FMAP_74_13);
			MULT_14(73)<=signed(DIN_14_7)*signed(FMAP_74_14);
			MULT_15(73)<=signed(DIN_15_7)*signed(FMAP_74_15);
			MULT_16(73)<=signed(DIN_16_7)*signed(FMAP_74_16);
			MULT_17(73)<=signed(DIN_17_7)*signed(FMAP_74_17);
			MULT_18(73)<=signed(DIN_18_7)*signed(FMAP_74_18);
			MULT_19(73)<=signed(DIN_19_7)*signed(FMAP_74_19);
			MULT_20(73)<=signed(DIN_20_7)*signed(FMAP_74_20);
			MULT_21(73)<=signed(DIN_21_7)*signed(FMAP_74_21);
			MULT_22(73)<=signed(DIN_22_7)*signed(FMAP_74_22);
			MULT_23(73)<=signed(DIN_23_7)*signed(FMAP_74_23);
			MULT_24(73)<=signed(DIN_24_7)*signed(FMAP_74_24);
			MULT_25(73)<=signed(DIN_25_7)*signed(FMAP_74_25);
			MULT_26(73)<=signed(DIN_26_7)*signed(FMAP_74_26);
			MULT_27(73)<=signed(DIN_27_7)*signed(FMAP_74_27);
			MULT_28(73)<=signed(DIN_28_7)*signed(FMAP_74_28);
			MULT_29(73)<=signed(DIN_29_7)*signed(FMAP_74_29);
			MULT_30(73)<=signed(DIN_30_7)*signed(FMAP_74_30);
			MULT_31(73)<=signed(DIN_31_7)*signed(FMAP_74_31);
			MULT_32(73)<=signed(DIN_32_7)*signed(FMAP_74_32);
			MULT_33(73)<=signed(DIN_33_7)*signed(FMAP_74_33);
			MULT_34(73)<=signed(DIN_34_7)*signed(FMAP_74_34);
			MULT_35(73)<=signed(DIN_35_7)*signed(FMAP_74_35);
			MULT_36(73)<=signed(DIN_36_7)*signed(FMAP_74_36);
			MULT_37(73)<=signed(DIN_37_7)*signed(FMAP_74_37);
			MULT_38(73)<=signed(DIN_38_7)*signed(FMAP_74_38);
			MULT_39(73)<=signed(DIN_39_7)*signed(FMAP_74_39);
			MULT_40(73)<=signed(DIN_40_7)*signed(FMAP_74_40);
			MULT_41(73)<=signed(DIN_41_7)*signed(FMAP_74_41);
			MULT_42(73)<=signed(DIN_42_7)*signed(FMAP_74_42);
			MULT_43(73)<=signed(DIN_43_7)*signed(FMAP_74_43);
			MULT_44(73)<=signed(DIN_44_7)*signed(FMAP_74_44);
			MULT_45(73)<=signed(DIN_45_7)*signed(FMAP_74_45);
			MULT_46(73)<=signed(DIN_46_7)*signed(FMAP_74_46);
			MULT_47(73)<=signed(DIN_47_7)*signed(FMAP_74_47);
			MULT_48(73)<=signed(DIN_48_7)*signed(FMAP_74_48);
			MULT_49(73)<=signed(DIN_49_7)*signed(FMAP_74_49);
			MULT_50(73)<=signed(DIN_50_7)*signed(FMAP_74_50);
			MULT_51(73)<=signed(DIN_51_7)*signed(FMAP_74_51);
			MULT_52(73)<=signed(DIN_52_7)*signed(FMAP_74_52);
			MULT_53(73)<=signed(DIN_53_7)*signed(FMAP_74_53);
			MULT_54(73)<=signed(DIN_54_7)*signed(FMAP_74_54);
			MULT_55(73)<=signed(DIN_55_7)*signed(FMAP_74_55);
			MULT_56(73)<=signed(DIN_56_7)*signed(FMAP_74_56);
			MULT_57(73)<=signed(DIN_57_7)*signed(FMAP_74_57);
			MULT_58(73)<=signed(DIN_58_7)*signed(FMAP_74_58);
			MULT_59(73)<=signed(DIN_59_7)*signed(FMAP_74_59);
			MULT_60(73)<=signed(DIN_60_7)*signed(FMAP_74_60);
			MULT_61(73)<=signed(DIN_61_7)*signed(FMAP_74_61);
			MULT_62(73)<=signed(DIN_62_7)*signed(FMAP_74_62);
			MULT_63(73)<=signed(DIN_63_7)*signed(FMAP_74_63);
			MULT_64(73)<=signed(DIN_64_7)*signed(FMAP_74_64);
			MULT_65(73)<=signed(DIN_65_7)*signed(FMAP_74_65);
			MULT_66(73)<=signed(DIN_66_7)*signed(FMAP_74_66);
			MULT_67(73)<=signed(DIN_67_7)*signed(FMAP_74_67);
			MULT_68(73)<=signed(DIN_68_7)*signed(FMAP_74_68);
			MULT_69(73)<=signed(DIN_69_7)*signed(FMAP_74_69);
			MULT_70(73)<=signed(DIN_70_7)*signed(FMAP_74_70);
			MULT_71(73)<=signed(DIN_71_7)*signed(FMAP_74_71);
			MULT_72(73)<=signed(DIN_72_7)*signed(FMAP_74_72);
			MULT_73(73)<=signed(DIN_73_7)*signed(FMAP_74_73);
			MULT_74(73)<=signed(DIN_74_7)*signed(FMAP_74_74);
			MULT_75(73)<=signed(DIN_75_7)*signed(FMAP_74_75);
			MULT_76(73)<=signed(DIN_76_7)*signed(FMAP_74_76);
			MULT_77(73)<=signed(DIN_77_7)*signed(FMAP_74_77);
			MULT_78(73)<=signed(DIN_78_7)*signed(FMAP_74_78);
			MULT_79(73)<=signed(DIN_79_7)*signed(FMAP_74_79);
			MULT_80(73)<=signed(DIN_80_7)*signed(FMAP_74_80);
			MULT_81(73)<=signed(DIN_81_7)*signed(FMAP_74_81);
			MULT_82(73)<=signed(DIN_82_7)*signed(FMAP_74_82);
			MULT_83(73)<=signed(DIN_83_7)*signed(FMAP_74_83);
			MULT_84(73)<=signed(DIN_84_7)*signed(FMAP_74_84);
			MULT_85(73)<=signed(DIN_85_7)*signed(FMAP_74_85);
			MULT_86(73)<=signed(DIN_86_7)*signed(FMAP_74_86);
			MULT_87(73)<=signed(DIN_87_7)*signed(FMAP_74_87);
			MULT_88(73)<=signed(DIN_88_7)*signed(FMAP_74_88);
			MULT_89(73)<=signed(DIN_89_7)*signed(FMAP_74_89);
			MULT_90(73)<=signed(DIN_90_7)*signed(FMAP_74_90);
			MULT_91(73)<=signed(DIN_91_7)*signed(FMAP_74_91);
			MULT_92(73)<=signed(DIN_92_7)*signed(FMAP_74_92);
			MULT_93(73)<=signed(DIN_93_7)*signed(FMAP_74_93);
			MULT_94(73)<=signed(DIN_94_7)*signed(FMAP_74_94);
			MULT_95(73)<=signed(DIN_95_7)*signed(FMAP_74_95);
			MULT_96(73)<=signed(DIN_96_7)*signed(FMAP_74_96);
			MULT_97(73)<=signed(DIN_97_7)*signed(FMAP_74_97);
			MULT_98(73)<=signed(DIN_98_7)*signed(FMAP_74_98);
			MULT_99(73)<=signed(DIN_99_7)*signed(FMAP_74_99);
			MULT_100(73)<=signed(DIN_100_7)*signed(FMAP_74_100);
			MULT_101(73)<=signed(DIN_101_7)*signed(FMAP_74_101);
			MULT_102(73)<=signed(DIN_102_7)*signed(FMAP_74_102);
			MULT_103(73)<=signed(DIN_103_7)*signed(FMAP_74_103);
			MULT_104(73)<=signed(DIN_104_7)*signed(FMAP_74_104);
			MULT_105(73)<=signed(DIN_105_7)*signed(FMAP_74_105);
			MULT_106(73)<=signed(DIN_106_7)*signed(FMAP_74_106);
			MULT_107(73)<=signed(DIN_107_7)*signed(FMAP_74_107);
			MULT_108(73)<=signed(DIN_108_7)*signed(FMAP_74_108);
			MULT_109(73)<=signed(DIN_109_7)*signed(FMAP_74_109);
			MULT_110(73)<=signed(DIN_110_7)*signed(FMAP_74_110);
			MULT_111(73)<=signed(DIN_111_7)*signed(FMAP_74_111);
			MULT_112(73)<=signed(DIN_112_7)*signed(FMAP_74_112);
			MULT_113(73)<=signed(DIN_113_7)*signed(FMAP_74_113);
			MULT_114(73)<=signed(DIN_114_7)*signed(FMAP_74_114);
			MULT_115(73)<=signed(DIN_115_7)*signed(FMAP_74_115);
			MULT_116(73)<=signed(DIN_116_7)*signed(FMAP_74_116);
			MULT_117(73)<=signed(DIN_117_7)*signed(FMAP_74_117);
			MULT_118(73)<=signed(DIN_118_7)*signed(FMAP_74_118);
			MULT_119(73)<=signed(DIN_119_7)*signed(FMAP_74_119);
			MULT_120(73)<=signed(DIN_120_7)*signed(FMAP_74_120);

			MULT_1(74)<=signed(DIN_1_7)*signed(FMAP_75_1);
			MULT_2(74)<=signed(DIN_2_7)*signed(FMAP_75_2);
			MULT_3(74)<=signed(DIN_3_7)*signed(FMAP_75_3);
			MULT_4(74)<=signed(DIN_4_7)*signed(FMAP_75_4);
			MULT_5(74)<=signed(DIN_5_7)*signed(FMAP_75_5);
			MULT_6(74)<=signed(DIN_6_7)*signed(FMAP_75_6);
			MULT_7(74)<=signed(DIN_7_7)*signed(FMAP_75_7);
			MULT_8(74)<=signed(DIN_8_7)*signed(FMAP_75_8);
			MULT_9(74)<=signed(DIN_9_7)*signed(FMAP_75_9);
			MULT_10(74)<=signed(DIN_10_7)*signed(FMAP_75_10);
			MULT_11(74)<=signed(DIN_11_7)*signed(FMAP_75_11);
			MULT_12(74)<=signed(DIN_12_7)*signed(FMAP_75_12);
			MULT_13(74)<=signed(DIN_13_7)*signed(FMAP_75_13);
			MULT_14(74)<=signed(DIN_14_7)*signed(FMAP_75_14);
			MULT_15(74)<=signed(DIN_15_7)*signed(FMAP_75_15);
			MULT_16(74)<=signed(DIN_16_7)*signed(FMAP_75_16);
			MULT_17(74)<=signed(DIN_17_7)*signed(FMAP_75_17);
			MULT_18(74)<=signed(DIN_18_7)*signed(FMAP_75_18);
			MULT_19(74)<=signed(DIN_19_7)*signed(FMAP_75_19);
			MULT_20(74)<=signed(DIN_20_7)*signed(FMAP_75_20);
			MULT_21(74)<=signed(DIN_21_7)*signed(FMAP_75_21);
			MULT_22(74)<=signed(DIN_22_7)*signed(FMAP_75_22);
			MULT_23(74)<=signed(DIN_23_7)*signed(FMAP_75_23);
			MULT_24(74)<=signed(DIN_24_7)*signed(FMAP_75_24);
			MULT_25(74)<=signed(DIN_25_7)*signed(FMAP_75_25);
			MULT_26(74)<=signed(DIN_26_7)*signed(FMAP_75_26);
			MULT_27(74)<=signed(DIN_27_7)*signed(FMAP_75_27);
			MULT_28(74)<=signed(DIN_28_7)*signed(FMAP_75_28);
			MULT_29(74)<=signed(DIN_29_7)*signed(FMAP_75_29);
			MULT_30(74)<=signed(DIN_30_7)*signed(FMAP_75_30);
			MULT_31(74)<=signed(DIN_31_7)*signed(FMAP_75_31);
			MULT_32(74)<=signed(DIN_32_7)*signed(FMAP_75_32);
			MULT_33(74)<=signed(DIN_33_7)*signed(FMAP_75_33);
			MULT_34(74)<=signed(DIN_34_7)*signed(FMAP_75_34);
			MULT_35(74)<=signed(DIN_35_7)*signed(FMAP_75_35);
			MULT_36(74)<=signed(DIN_36_7)*signed(FMAP_75_36);
			MULT_37(74)<=signed(DIN_37_7)*signed(FMAP_75_37);
			MULT_38(74)<=signed(DIN_38_7)*signed(FMAP_75_38);
			MULT_39(74)<=signed(DIN_39_7)*signed(FMAP_75_39);
			MULT_40(74)<=signed(DIN_40_7)*signed(FMAP_75_40);
			MULT_41(74)<=signed(DIN_41_7)*signed(FMAP_75_41);
			MULT_42(74)<=signed(DIN_42_7)*signed(FMAP_75_42);
			MULT_43(74)<=signed(DIN_43_7)*signed(FMAP_75_43);
			MULT_44(74)<=signed(DIN_44_7)*signed(FMAP_75_44);
			MULT_45(74)<=signed(DIN_45_7)*signed(FMAP_75_45);
			MULT_46(74)<=signed(DIN_46_7)*signed(FMAP_75_46);
			MULT_47(74)<=signed(DIN_47_7)*signed(FMAP_75_47);
			MULT_48(74)<=signed(DIN_48_7)*signed(FMAP_75_48);
			MULT_49(74)<=signed(DIN_49_7)*signed(FMAP_75_49);
			MULT_50(74)<=signed(DIN_50_7)*signed(FMAP_75_50);
			MULT_51(74)<=signed(DIN_51_7)*signed(FMAP_75_51);
			MULT_52(74)<=signed(DIN_52_7)*signed(FMAP_75_52);
			MULT_53(74)<=signed(DIN_53_7)*signed(FMAP_75_53);
			MULT_54(74)<=signed(DIN_54_7)*signed(FMAP_75_54);
			MULT_55(74)<=signed(DIN_55_7)*signed(FMAP_75_55);
			MULT_56(74)<=signed(DIN_56_7)*signed(FMAP_75_56);
			MULT_57(74)<=signed(DIN_57_7)*signed(FMAP_75_57);
			MULT_58(74)<=signed(DIN_58_7)*signed(FMAP_75_58);
			MULT_59(74)<=signed(DIN_59_7)*signed(FMAP_75_59);
			MULT_60(74)<=signed(DIN_60_7)*signed(FMAP_75_60);
			MULT_61(74)<=signed(DIN_61_7)*signed(FMAP_75_61);
			MULT_62(74)<=signed(DIN_62_7)*signed(FMAP_75_62);
			MULT_63(74)<=signed(DIN_63_7)*signed(FMAP_75_63);
			MULT_64(74)<=signed(DIN_64_7)*signed(FMAP_75_64);
			MULT_65(74)<=signed(DIN_65_7)*signed(FMAP_75_65);
			MULT_66(74)<=signed(DIN_66_7)*signed(FMAP_75_66);
			MULT_67(74)<=signed(DIN_67_7)*signed(FMAP_75_67);
			MULT_68(74)<=signed(DIN_68_7)*signed(FMAP_75_68);
			MULT_69(74)<=signed(DIN_69_7)*signed(FMAP_75_69);
			MULT_70(74)<=signed(DIN_70_7)*signed(FMAP_75_70);
			MULT_71(74)<=signed(DIN_71_7)*signed(FMAP_75_71);
			MULT_72(74)<=signed(DIN_72_7)*signed(FMAP_75_72);
			MULT_73(74)<=signed(DIN_73_7)*signed(FMAP_75_73);
			MULT_74(74)<=signed(DIN_74_7)*signed(FMAP_75_74);
			MULT_75(74)<=signed(DIN_75_7)*signed(FMAP_75_75);
			MULT_76(74)<=signed(DIN_76_7)*signed(FMAP_75_76);
			MULT_77(74)<=signed(DIN_77_7)*signed(FMAP_75_77);
			MULT_78(74)<=signed(DIN_78_7)*signed(FMAP_75_78);
			MULT_79(74)<=signed(DIN_79_7)*signed(FMAP_75_79);
			MULT_80(74)<=signed(DIN_80_7)*signed(FMAP_75_80);
			MULT_81(74)<=signed(DIN_81_7)*signed(FMAP_75_81);
			MULT_82(74)<=signed(DIN_82_7)*signed(FMAP_75_82);
			MULT_83(74)<=signed(DIN_83_7)*signed(FMAP_75_83);
			MULT_84(74)<=signed(DIN_84_7)*signed(FMAP_75_84);
			MULT_85(74)<=signed(DIN_85_7)*signed(FMAP_75_85);
			MULT_86(74)<=signed(DIN_86_7)*signed(FMAP_75_86);
			MULT_87(74)<=signed(DIN_87_7)*signed(FMAP_75_87);
			MULT_88(74)<=signed(DIN_88_7)*signed(FMAP_75_88);
			MULT_89(74)<=signed(DIN_89_7)*signed(FMAP_75_89);
			MULT_90(74)<=signed(DIN_90_7)*signed(FMAP_75_90);
			MULT_91(74)<=signed(DIN_91_7)*signed(FMAP_75_91);
			MULT_92(74)<=signed(DIN_92_7)*signed(FMAP_75_92);
			MULT_93(74)<=signed(DIN_93_7)*signed(FMAP_75_93);
			MULT_94(74)<=signed(DIN_94_7)*signed(FMAP_75_94);
			MULT_95(74)<=signed(DIN_95_7)*signed(FMAP_75_95);
			MULT_96(74)<=signed(DIN_96_7)*signed(FMAP_75_96);
			MULT_97(74)<=signed(DIN_97_7)*signed(FMAP_75_97);
			MULT_98(74)<=signed(DIN_98_7)*signed(FMAP_75_98);
			MULT_99(74)<=signed(DIN_99_7)*signed(FMAP_75_99);
			MULT_100(74)<=signed(DIN_100_7)*signed(FMAP_75_100);
			MULT_101(74)<=signed(DIN_101_7)*signed(FMAP_75_101);
			MULT_102(74)<=signed(DIN_102_7)*signed(FMAP_75_102);
			MULT_103(74)<=signed(DIN_103_7)*signed(FMAP_75_103);
			MULT_104(74)<=signed(DIN_104_7)*signed(FMAP_75_104);
			MULT_105(74)<=signed(DIN_105_7)*signed(FMAP_75_105);
			MULT_106(74)<=signed(DIN_106_7)*signed(FMAP_75_106);
			MULT_107(74)<=signed(DIN_107_7)*signed(FMAP_75_107);
			MULT_108(74)<=signed(DIN_108_7)*signed(FMAP_75_108);
			MULT_109(74)<=signed(DIN_109_7)*signed(FMAP_75_109);
			MULT_110(74)<=signed(DIN_110_7)*signed(FMAP_75_110);
			MULT_111(74)<=signed(DIN_111_7)*signed(FMAP_75_111);
			MULT_112(74)<=signed(DIN_112_7)*signed(FMAP_75_112);
			MULT_113(74)<=signed(DIN_113_7)*signed(FMAP_75_113);
			MULT_114(74)<=signed(DIN_114_7)*signed(FMAP_75_114);
			MULT_115(74)<=signed(DIN_115_7)*signed(FMAP_75_115);
			MULT_116(74)<=signed(DIN_116_7)*signed(FMAP_75_116);
			MULT_117(74)<=signed(DIN_117_7)*signed(FMAP_75_117);
			MULT_118(74)<=signed(DIN_118_7)*signed(FMAP_75_118);
			MULT_119(74)<=signed(DIN_119_7)*signed(FMAP_75_119);
			MULT_120(74)<=signed(DIN_120_7)*signed(FMAP_75_120);

			MULT_1(75)<=signed(DIN_1_7)*signed(FMAP_76_1);
			MULT_2(75)<=signed(DIN_2_7)*signed(FMAP_76_2);
			MULT_3(75)<=signed(DIN_3_7)*signed(FMAP_76_3);
			MULT_4(75)<=signed(DIN_4_7)*signed(FMAP_76_4);
			MULT_5(75)<=signed(DIN_5_7)*signed(FMAP_76_5);
			MULT_6(75)<=signed(DIN_6_7)*signed(FMAP_76_6);
			MULT_7(75)<=signed(DIN_7_7)*signed(FMAP_76_7);
			MULT_8(75)<=signed(DIN_8_7)*signed(FMAP_76_8);
			MULT_9(75)<=signed(DIN_9_7)*signed(FMAP_76_9);
			MULT_10(75)<=signed(DIN_10_7)*signed(FMAP_76_10);
			MULT_11(75)<=signed(DIN_11_7)*signed(FMAP_76_11);
			MULT_12(75)<=signed(DIN_12_7)*signed(FMAP_76_12);
			MULT_13(75)<=signed(DIN_13_7)*signed(FMAP_76_13);
			MULT_14(75)<=signed(DIN_14_7)*signed(FMAP_76_14);
			MULT_15(75)<=signed(DIN_15_7)*signed(FMAP_76_15);
			MULT_16(75)<=signed(DIN_16_7)*signed(FMAP_76_16);
			MULT_17(75)<=signed(DIN_17_7)*signed(FMAP_76_17);
			MULT_18(75)<=signed(DIN_18_7)*signed(FMAP_76_18);
			MULT_19(75)<=signed(DIN_19_7)*signed(FMAP_76_19);
			MULT_20(75)<=signed(DIN_20_7)*signed(FMAP_76_20);
			MULT_21(75)<=signed(DIN_21_7)*signed(FMAP_76_21);
			MULT_22(75)<=signed(DIN_22_7)*signed(FMAP_76_22);
			MULT_23(75)<=signed(DIN_23_7)*signed(FMAP_76_23);
			MULT_24(75)<=signed(DIN_24_7)*signed(FMAP_76_24);
			MULT_25(75)<=signed(DIN_25_7)*signed(FMAP_76_25);
			MULT_26(75)<=signed(DIN_26_7)*signed(FMAP_76_26);
			MULT_27(75)<=signed(DIN_27_7)*signed(FMAP_76_27);
			MULT_28(75)<=signed(DIN_28_7)*signed(FMAP_76_28);
			MULT_29(75)<=signed(DIN_29_7)*signed(FMAP_76_29);
			MULT_30(75)<=signed(DIN_30_7)*signed(FMAP_76_30);
			MULT_31(75)<=signed(DIN_31_7)*signed(FMAP_76_31);
			MULT_32(75)<=signed(DIN_32_7)*signed(FMAP_76_32);
			MULT_33(75)<=signed(DIN_33_7)*signed(FMAP_76_33);
			MULT_34(75)<=signed(DIN_34_7)*signed(FMAP_76_34);
			MULT_35(75)<=signed(DIN_35_7)*signed(FMAP_76_35);
			MULT_36(75)<=signed(DIN_36_7)*signed(FMAP_76_36);
			MULT_37(75)<=signed(DIN_37_7)*signed(FMAP_76_37);
			MULT_38(75)<=signed(DIN_38_7)*signed(FMAP_76_38);
			MULT_39(75)<=signed(DIN_39_7)*signed(FMAP_76_39);
			MULT_40(75)<=signed(DIN_40_7)*signed(FMAP_76_40);
			MULT_41(75)<=signed(DIN_41_7)*signed(FMAP_76_41);
			MULT_42(75)<=signed(DIN_42_7)*signed(FMAP_76_42);
			MULT_43(75)<=signed(DIN_43_7)*signed(FMAP_76_43);
			MULT_44(75)<=signed(DIN_44_7)*signed(FMAP_76_44);
			MULT_45(75)<=signed(DIN_45_7)*signed(FMAP_76_45);
			MULT_46(75)<=signed(DIN_46_7)*signed(FMAP_76_46);
			MULT_47(75)<=signed(DIN_47_7)*signed(FMAP_76_47);
			MULT_48(75)<=signed(DIN_48_7)*signed(FMAP_76_48);
			MULT_49(75)<=signed(DIN_49_7)*signed(FMAP_76_49);
			MULT_50(75)<=signed(DIN_50_7)*signed(FMAP_76_50);
			MULT_51(75)<=signed(DIN_51_7)*signed(FMAP_76_51);
			MULT_52(75)<=signed(DIN_52_7)*signed(FMAP_76_52);
			MULT_53(75)<=signed(DIN_53_7)*signed(FMAP_76_53);
			MULT_54(75)<=signed(DIN_54_7)*signed(FMAP_76_54);
			MULT_55(75)<=signed(DIN_55_7)*signed(FMAP_76_55);
			MULT_56(75)<=signed(DIN_56_7)*signed(FMAP_76_56);
			MULT_57(75)<=signed(DIN_57_7)*signed(FMAP_76_57);
			MULT_58(75)<=signed(DIN_58_7)*signed(FMAP_76_58);
			MULT_59(75)<=signed(DIN_59_7)*signed(FMAP_76_59);
			MULT_60(75)<=signed(DIN_60_7)*signed(FMAP_76_60);
			MULT_61(75)<=signed(DIN_61_7)*signed(FMAP_76_61);
			MULT_62(75)<=signed(DIN_62_7)*signed(FMAP_76_62);
			MULT_63(75)<=signed(DIN_63_7)*signed(FMAP_76_63);
			MULT_64(75)<=signed(DIN_64_7)*signed(FMAP_76_64);
			MULT_65(75)<=signed(DIN_65_7)*signed(FMAP_76_65);
			MULT_66(75)<=signed(DIN_66_7)*signed(FMAP_76_66);
			MULT_67(75)<=signed(DIN_67_7)*signed(FMAP_76_67);
			MULT_68(75)<=signed(DIN_68_7)*signed(FMAP_76_68);
			MULT_69(75)<=signed(DIN_69_7)*signed(FMAP_76_69);
			MULT_70(75)<=signed(DIN_70_7)*signed(FMAP_76_70);
			MULT_71(75)<=signed(DIN_71_7)*signed(FMAP_76_71);
			MULT_72(75)<=signed(DIN_72_7)*signed(FMAP_76_72);
			MULT_73(75)<=signed(DIN_73_7)*signed(FMAP_76_73);
			MULT_74(75)<=signed(DIN_74_7)*signed(FMAP_76_74);
			MULT_75(75)<=signed(DIN_75_7)*signed(FMAP_76_75);
			MULT_76(75)<=signed(DIN_76_7)*signed(FMAP_76_76);
			MULT_77(75)<=signed(DIN_77_7)*signed(FMAP_76_77);
			MULT_78(75)<=signed(DIN_78_7)*signed(FMAP_76_78);
			MULT_79(75)<=signed(DIN_79_7)*signed(FMAP_76_79);
			MULT_80(75)<=signed(DIN_80_7)*signed(FMAP_76_80);
			MULT_81(75)<=signed(DIN_81_7)*signed(FMAP_76_81);
			MULT_82(75)<=signed(DIN_82_7)*signed(FMAP_76_82);
			MULT_83(75)<=signed(DIN_83_7)*signed(FMAP_76_83);
			MULT_84(75)<=signed(DIN_84_7)*signed(FMAP_76_84);
			MULT_85(75)<=signed(DIN_85_7)*signed(FMAP_76_85);
			MULT_86(75)<=signed(DIN_86_7)*signed(FMAP_76_86);
			MULT_87(75)<=signed(DIN_87_7)*signed(FMAP_76_87);
			MULT_88(75)<=signed(DIN_88_7)*signed(FMAP_76_88);
			MULT_89(75)<=signed(DIN_89_7)*signed(FMAP_76_89);
			MULT_90(75)<=signed(DIN_90_7)*signed(FMAP_76_90);
			MULT_91(75)<=signed(DIN_91_7)*signed(FMAP_76_91);
			MULT_92(75)<=signed(DIN_92_7)*signed(FMAP_76_92);
			MULT_93(75)<=signed(DIN_93_7)*signed(FMAP_76_93);
			MULT_94(75)<=signed(DIN_94_7)*signed(FMAP_76_94);
			MULT_95(75)<=signed(DIN_95_7)*signed(FMAP_76_95);
			MULT_96(75)<=signed(DIN_96_7)*signed(FMAP_76_96);
			MULT_97(75)<=signed(DIN_97_7)*signed(FMAP_76_97);
			MULT_98(75)<=signed(DIN_98_7)*signed(FMAP_76_98);
			MULT_99(75)<=signed(DIN_99_7)*signed(FMAP_76_99);
			MULT_100(75)<=signed(DIN_100_7)*signed(FMAP_76_100);
			MULT_101(75)<=signed(DIN_101_7)*signed(FMAP_76_101);
			MULT_102(75)<=signed(DIN_102_7)*signed(FMAP_76_102);
			MULT_103(75)<=signed(DIN_103_7)*signed(FMAP_76_103);
			MULT_104(75)<=signed(DIN_104_7)*signed(FMAP_76_104);
			MULT_105(75)<=signed(DIN_105_7)*signed(FMAP_76_105);
			MULT_106(75)<=signed(DIN_106_7)*signed(FMAP_76_106);
			MULT_107(75)<=signed(DIN_107_7)*signed(FMAP_76_107);
			MULT_108(75)<=signed(DIN_108_7)*signed(FMAP_76_108);
			MULT_109(75)<=signed(DIN_109_7)*signed(FMAP_76_109);
			MULT_110(75)<=signed(DIN_110_7)*signed(FMAP_76_110);
			MULT_111(75)<=signed(DIN_111_7)*signed(FMAP_76_111);
			MULT_112(75)<=signed(DIN_112_7)*signed(FMAP_76_112);
			MULT_113(75)<=signed(DIN_113_7)*signed(FMAP_76_113);
			MULT_114(75)<=signed(DIN_114_7)*signed(FMAP_76_114);
			MULT_115(75)<=signed(DIN_115_7)*signed(FMAP_76_115);
			MULT_116(75)<=signed(DIN_116_7)*signed(FMAP_76_116);
			MULT_117(75)<=signed(DIN_117_7)*signed(FMAP_76_117);
			MULT_118(75)<=signed(DIN_118_7)*signed(FMAP_76_118);
			MULT_119(75)<=signed(DIN_119_7)*signed(FMAP_76_119);
			MULT_120(75)<=signed(DIN_120_7)*signed(FMAP_76_120);

			MULT_1(76)<=signed(DIN_1_7)*signed(FMAP_77_1);
			MULT_2(76)<=signed(DIN_2_7)*signed(FMAP_77_2);
			MULT_3(76)<=signed(DIN_3_7)*signed(FMAP_77_3);
			MULT_4(76)<=signed(DIN_4_7)*signed(FMAP_77_4);
			MULT_5(76)<=signed(DIN_5_7)*signed(FMAP_77_5);
			MULT_6(76)<=signed(DIN_6_7)*signed(FMAP_77_6);
			MULT_7(76)<=signed(DIN_7_7)*signed(FMAP_77_7);
			MULT_8(76)<=signed(DIN_8_7)*signed(FMAP_77_8);
			MULT_9(76)<=signed(DIN_9_7)*signed(FMAP_77_9);
			MULT_10(76)<=signed(DIN_10_7)*signed(FMAP_77_10);
			MULT_11(76)<=signed(DIN_11_7)*signed(FMAP_77_11);
			MULT_12(76)<=signed(DIN_12_7)*signed(FMAP_77_12);
			MULT_13(76)<=signed(DIN_13_7)*signed(FMAP_77_13);
			MULT_14(76)<=signed(DIN_14_7)*signed(FMAP_77_14);
			MULT_15(76)<=signed(DIN_15_7)*signed(FMAP_77_15);
			MULT_16(76)<=signed(DIN_16_7)*signed(FMAP_77_16);
			MULT_17(76)<=signed(DIN_17_7)*signed(FMAP_77_17);
			MULT_18(76)<=signed(DIN_18_7)*signed(FMAP_77_18);
			MULT_19(76)<=signed(DIN_19_7)*signed(FMAP_77_19);
			MULT_20(76)<=signed(DIN_20_7)*signed(FMAP_77_20);
			MULT_21(76)<=signed(DIN_21_7)*signed(FMAP_77_21);
			MULT_22(76)<=signed(DIN_22_7)*signed(FMAP_77_22);
			MULT_23(76)<=signed(DIN_23_7)*signed(FMAP_77_23);
			MULT_24(76)<=signed(DIN_24_7)*signed(FMAP_77_24);
			MULT_25(76)<=signed(DIN_25_7)*signed(FMAP_77_25);
			MULT_26(76)<=signed(DIN_26_7)*signed(FMAP_77_26);
			MULT_27(76)<=signed(DIN_27_7)*signed(FMAP_77_27);
			MULT_28(76)<=signed(DIN_28_7)*signed(FMAP_77_28);
			MULT_29(76)<=signed(DIN_29_7)*signed(FMAP_77_29);
			MULT_30(76)<=signed(DIN_30_7)*signed(FMAP_77_30);
			MULT_31(76)<=signed(DIN_31_7)*signed(FMAP_77_31);
			MULT_32(76)<=signed(DIN_32_7)*signed(FMAP_77_32);
			MULT_33(76)<=signed(DIN_33_7)*signed(FMAP_77_33);
			MULT_34(76)<=signed(DIN_34_7)*signed(FMAP_77_34);
			MULT_35(76)<=signed(DIN_35_7)*signed(FMAP_77_35);
			MULT_36(76)<=signed(DIN_36_7)*signed(FMAP_77_36);
			MULT_37(76)<=signed(DIN_37_7)*signed(FMAP_77_37);
			MULT_38(76)<=signed(DIN_38_7)*signed(FMAP_77_38);
			MULT_39(76)<=signed(DIN_39_7)*signed(FMAP_77_39);
			MULT_40(76)<=signed(DIN_40_7)*signed(FMAP_77_40);
			MULT_41(76)<=signed(DIN_41_7)*signed(FMAP_77_41);
			MULT_42(76)<=signed(DIN_42_7)*signed(FMAP_77_42);
			MULT_43(76)<=signed(DIN_43_7)*signed(FMAP_77_43);
			MULT_44(76)<=signed(DIN_44_7)*signed(FMAP_77_44);
			MULT_45(76)<=signed(DIN_45_7)*signed(FMAP_77_45);
			MULT_46(76)<=signed(DIN_46_7)*signed(FMAP_77_46);
			MULT_47(76)<=signed(DIN_47_7)*signed(FMAP_77_47);
			MULT_48(76)<=signed(DIN_48_7)*signed(FMAP_77_48);
			MULT_49(76)<=signed(DIN_49_7)*signed(FMAP_77_49);
			MULT_50(76)<=signed(DIN_50_7)*signed(FMAP_77_50);
			MULT_51(76)<=signed(DIN_51_7)*signed(FMAP_77_51);
			MULT_52(76)<=signed(DIN_52_7)*signed(FMAP_77_52);
			MULT_53(76)<=signed(DIN_53_7)*signed(FMAP_77_53);
			MULT_54(76)<=signed(DIN_54_7)*signed(FMAP_77_54);
			MULT_55(76)<=signed(DIN_55_7)*signed(FMAP_77_55);
			MULT_56(76)<=signed(DIN_56_7)*signed(FMAP_77_56);
			MULT_57(76)<=signed(DIN_57_7)*signed(FMAP_77_57);
			MULT_58(76)<=signed(DIN_58_7)*signed(FMAP_77_58);
			MULT_59(76)<=signed(DIN_59_7)*signed(FMAP_77_59);
			MULT_60(76)<=signed(DIN_60_7)*signed(FMAP_77_60);
			MULT_61(76)<=signed(DIN_61_7)*signed(FMAP_77_61);
			MULT_62(76)<=signed(DIN_62_7)*signed(FMAP_77_62);
			MULT_63(76)<=signed(DIN_63_7)*signed(FMAP_77_63);
			MULT_64(76)<=signed(DIN_64_7)*signed(FMAP_77_64);
			MULT_65(76)<=signed(DIN_65_7)*signed(FMAP_77_65);
			MULT_66(76)<=signed(DIN_66_7)*signed(FMAP_77_66);
			MULT_67(76)<=signed(DIN_67_7)*signed(FMAP_77_67);
			MULT_68(76)<=signed(DIN_68_7)*signed(FMAP_77_68);
			MULT_69(76)<=signed(DIN_69_7)*signed(FMAP_77_69);
			MULT_70(76)<=signed(DIN_70_7)*signed(FMAP_77_70);
			MULT_71(76)<=signed(DIN_71_7)*signed(FMAP_77_71);
			MULT_72(76)<=signed(DIN_72_7)*signed(FMAP_77_72);
			MULT_73(76)<=signed(DIN_73_7)*signed(FMAP_77_73);
			MULT_74(76)<=signed(DIN_74_7)*signed(FMAP_77_74);
			MULT_75(76)<=signed(DIN_75_7)*signed(FMAP_77_75);
			MULT_76(76)<=signed(DIN_76_7)*signed(FMAP_77_76);
			MULT_77(76)<=signed(DIN_77_7)*signed(FMAP_77_77);
			MULT_78(76)<=signed(DIN_78_7)*signed(FMAP_77_78);
			MULT_79(76)<=signed(DIN_79_7)*signed(FMAP_77_79);
			MULT_80(76)<=signed(DIN_80_7)*signed(FMAP_77_80);
			MULT_81(76)<=signed(DIN_81_7)*signed(FMAP_77_81);
			MULT_82(76)<=signed(DIN_82_7)*signed(FMAP_77_82);
			MULT_83(76)<=signed(DIN_83_7)*signed(FMAP_77_83);
			MULT_84(76)<=signed(DIN_84_7)*signed(FMAP_77_84);
			MULT_85(76)<=signed(DIN_85_7)*signed(FMAP_77_85);
			MULT_86(76)<=signed(DIN_86_7)*signed(FMAP_77_86);
			MULT_87(76)<=signed(DIN_87_7)*signed(FMAP_77_87);
			MULT_88(76)<=signed(DIN_88_7)*signed(FMAP_77_88);
			MULT_89(76)<=signed(DIN_89_7)*signed(FMAP_77_89);
			MULT_90(76)<=signed(DIN_90_7)*signed(FMAP_77_90);
			MULT_91(76)<=signed(DIN_91_7)*signed(FMAP_77_91);
			MULT_92(76)<=signed(DIN_92_7)*signed(FMAP_77_92);
			MULT_93(76)<=signed(DIN_93_7)*signed(FMAP_77_93);
			MULT_94(76)<=signed(DIN_94_7)*signed(FMAP_77_94);
			MULT_95(76)<=signed(DIN_95_7)*signed(FMAP_77_95);
			MULT_96(76)<=signed(DIN_96_7)*signed(FMAP_77_96);
			MULT_97(76)<=signed(DIN_97_7)*signed(FMAP_77_97);
			MULT_98(76)<=signed(DIN_98_7)*signed(FMAP_77_98);
			MULT_99(76)<=signed(DIN_99_7)*signed(FMAP_77_99);
			MULT_100(76)<=signed(DIN_100_7)*signed(FMAP_77_100);
			MULT_101(76)<=signed(DIN_101_7)*signed(FMAP_77_101);
			MULT_102(76)<=signed(DIN_102_7)*signed(FMAP_77_102);
			MULT_103(76)<=signed(DIN_103_7)*signed(FMAP_77_103);
			MULT_104(76)<=signed(DIN_104_7)*signed(FMAP_77_104);
			MULT_105(76)<=signed(DIN_105_7)*signed(FMAP_77_105);
			MULT_106(76)<=signed(DIN_106_7)*signed(FMAP_77_106);
			MULT_107(76)<=signed(DIN_107_7)*signed(FMAP_77_107);
			MULT_108(76)<=signed(DIN_108_7)*signed(FMAP_77_108);
			MULT_109(76)<=signed(DIN_109_7)*signed(FMAP_77_109);
			MULT_110(76)<=signed(DIN_110_7)*signed(FMAP_77_110);
			MULT_111(76)<=signed(DIN_111_7)*signed(FMAP_77_111);
			MULT_112(76)<=signed(DIN_112_7)*signed(FMAP_77_112);
			MULT_113(76)<=signed(DIN_113_7)*signed(FMAP_77_113);
			MULT_114(76)<=signed(DIN_114_7)*signed(FMAP_77_114);
			MULT_115(76)<=signed(DIN_115_7)*signed(FMAP_77_115);
			MULT_116(76)<=signed(DIN_116_7)*signed(FMAP_77_116);
			MULT_117(76)<=signed(DIN_117_7)*signed(FMAP_77_117);
			MULT_118(76)<=signed(DIN_118_7)*signed(FMAP_77_118);
			MULT_119(76)<=signed(DIN_119_7)*signed(FMAP_77_119);
			MULT_120(76)<=signed(DIN_120_7)*signed(FMAP_77_120);

			MULT_1(77)<=signed(DIN_1_7)*signed(FMAP_78_1);
			MULT_2(77)<=signed(DIN_2_7)*signed(FMAP_78_2);
			MULT_3(77)<=signed(DIN_3_7)*signed(FMAP_78_3);
			MULT_4(77)<=signed(DIN_4_7)*signed(FMAP_78_4);
			MULT_5(77)<=signed(DIN_5_7)*signed(FMAP_78_5);
			MULT_6(77)<=signed(DIN_6_7)*signed(FMAP_78_6);
			MULT_7(77)<=signed(DIN_7_7)*signed(FMAP_78_7);
			MULT_8(77)<=signed(DIN_8_7)*signed(FMAP_78_8);
			MULT_9(77)<=signed(DIN_9_7)*signed(FMAP_78_9);
			MULT_10(77)<=signed(DIN_10_7)*signed(FMAP_78_10);
			MULT_11(77)<=signed(DIN_11_7)*signed(FMAP_78_11);
			MULT_12(77)<=signed(DIN_12_7)*signed(FMAP_78_12);
			MULT_13(77)<=signed(DIN_13_7)*signed(FMAP_78_13);
			MULT_14(77)<=signed(DIN_14_7)*signed(FMAP_78_14);
			MULT_15(77)<=signed(DIN_15_7)*signed(FMAP_78_15);
			MULT_16(77)<=signed(DIN_16_7)*signed(FMAP_78_16);
			MULT_17(77)<=signed(DIN_17_7)*signed(FMAP_78_17);
			MULT_18(77)<=signed(DIN_18_7)*signed(FMAP_78_18);
			MULT_19(77)<=signed(DIN_19_7)*signed(FMAP_78_19);
			MULT_20(77)<=signed(DIN_20_7)*signed(FMAP_78_20);
			MULT_21(77)<=signed(DIN_21_7)*signed(FMAP_78_21);
			MULT_22(77)<=signed(DIN_22_7)*signed(FMAP_78_22);
			MULT_23(77)<=signed(DIN_23_7)*signed(FMAP_78_23);
			MULT_24(77)<=signed(DIN_24_7)*signed(FMAP_78_24);
			MULT_25(77)<=signed(DIN_25_7)*signed(FMAP_78_25);
			MULT_26(77)<=signed(DIN_26_7)*signed(FMAP_78_26);
			MULT_27(77)<=signed(DIN_27_7)*signed(FMAP_78_27);
			MULT_28(77)<=signed(DIN_28_7)*signed(FMAP_78_28);
			MULT_29(77)<=signed(DIN_29_7)*signed(FMAP_78_29);
			MULT_30(77)<=signed(DIN_30_7)*signed(FMAP_78_30);
			MULT_31(77)<=signed(DIN_31_7)*signed(FMAP_78_31);
			MULT_32(77)<=signed(DIN_32_7)*signed(FMAP_78_32);
			MULT_33(77)<=signed(DIN_33_7)*signed(FMAP_78_33);
			MULT_34(77)<=signed(DIN_34_7)*signed(FMAP_78_34);
			MULT_35(77)<=signed(DIN_35_7)*signed(FMAP_78_35);
			MULT_36(77)<=signed(DIN_36_7)*signed(FMAP_78_36);
			MULT_37(77)<=signed(DIN_37_7)*signed(FMAP_78_37);
			MULT_38(77)<=signed(DIN_38_7)*signed(FMAP_78_38);
			MULT_39(77)<=signed(DIN_39_7)*signed(FMAP_78_39);
			MULT_40(77)<=signed(DIN_40_7)*signed(FMAP_78_40);
			MULT_41(77)<=signed(DIN_41_7)*signed(FMAP_78_41);
			MULT_42(77)<=signed(DIN_42_7)*signed(FMAP_78_42);
			MULT_43(77)<=signed(DIN_43_7)*signed(FMAP_78_43);
			MULT_44(77)<=signed(DIN_44_7)*signed(FMAP_78_44);
			MULT_45(77)<=signed(DIN_45_7)*signed(FMAP_78_45);
			MULT_46(77)<=signed(DIN_46_7)*signed(FMAP_78_46);
			MULT_47(77)<=signed(DIN_47_7)*signed(FMAP_78_47);
			MULT_48(77)<=signed(DIN_48_7)*signed(FMAP_78_48);
			MULT_49(77)<=signed(DIN_49_7)*signed(FMAP_78_49);
			MULT_50(77)<=signed(DIN_50_7)*signed(FMAP_78_50);
			MULT_51(77)<=signed(DIN_51_7)*signed(FMAP_78_51);
			MULT_52(77)<=signed(DIN_52_7)*signed(FMAP_78_52);
			MULT_53(77)<=signed(DIN_53_7)*signed(FMAP_78_53);
			MULT_54(77)<=signed(DIN_54_7)*signed(FMAP_78_54);
			MULT_55(77)<=signed(DIN_55_7)*signed(FMAP_78_55);
			MULT_56(77)<=signed(DIN_56_7)*signed(FMAP_78_56);
			MULT_57(77)<=signed(DIN_57_7)*signed(FMAP_78_57);
			MULT_58(77)<=signed(DIN_58_7)*signed(FMAP_78_58);
			MULT_59(77)<=signed(DIN_59_7)*signed(FMAP_78_59);
			MULT_60(77)<=signed(DIN_60_7)*signed(FMAP_78_60);
			MULT_61(77)<=signed(DIN_61_7)*signed(FMAP_78_61);
			MULT_62(77)<=signed(DIN_62_7)*signed(FMAP_78_62);
			MULT_63(77)<=signed(DIN_63_7)*signed(FMAP_78_63);
			MULT_64(77)<=signed(DIN_64_7)*signed(FMAP_78_64);
			MULT_65(77)<=signed(DIN_65_7)*signed(FMAP_78_65);
			MULT_66(77)<=signed(DIN_66_7)*signed(FMAP_78_66);
			MULT_67(77)<=signed(DIN_67_7)*signed(FMAP_78_67);
			MULT_68(77)<=signed(DIN_68_7)*signed(FMAP_78_68);
			MULT_69(77)<=signed(DIN_69_7)*signed(FMAP_78_69);
			MULT_70(77)<=signed(DIN_70_7)*signed(FMAP_78_70);
			MULT_71(77)<=signed(DIN_71_7)*signed(FMAP_78_71);
			MULT_72(77)<=signed(DIN_72_7)*signed(FMAP_78_72);
			MULT_73(77)<=signed(DIN_73_7)*signed(FMAP_78_73);
			MULT_74(77)<=signed(DIN_74_7)*signed(FMAP_78_74);
			MULT_75(77)<=signed(DIN_75_7)*signed(FMAP_78_75);
			MULT_76(77)<=signed(DIN_76_7)*signed(FMAP_78_76);
			MULT_77(77)<=signed(DIN_77_7)*signed(FMAP_78_77);
			MULT_78(77)<=signed(DIN_78_7)*signed(FMAP_78_78);
			MULT_79(77)<=signed(DIN_79_7)*signed(FMAP_78_79);
			MULT_80(77)<=signed(DIN_80_7)*signed(FMAP_78_80);
			MULT_81(77)<=signed(DIN_81_7)*signed(FMAP_78_81);
			MULT_82(77)<=signed(DIN_82_7)*signed(FMAP_78_82);
			MULT_83(77)<=signed(DIN_83_7)*signed(FMAP_78_83);
			MULT_84(77)<=signed(DIN_84_7)*signed(FMAP_78_84);
			MULT_85(77)<=signed(DIN_85_7)*signed(FMAP_78_85);
			MULT_86(77)<=signed(DIN_86_7)*signed(FMAP_78_86);
			MULT_87(77)<=signed(DIN_87_7)*signed(FMAP_78_87);
			MULT_88(77)<=signed(DIN_88_7)*signed(FMAP_78_88);
			MULT_89(77)<=signed(DIN_89_7)*signed(FMAP_78_89);
			MULT_90(77)<=signed(DIN_90_7)*signed(FMAP_78_90);
			MULT_91(77)<=signed(DIN_91_7)*signed(FMAP_78_91);
			MULT_92(77)<=signed(DIN_92_7)*signed(FMAP_78_92);
			MULT_93(77)<=signed(DIN_93_7)*signed(FMAP_78_93);
			MULT_94(77)<=signed(DIN_94_7)*signed(FMAP_78_94);
			MULT_95(77)<=signed(DIN_95_7)*signed(FMAP_78_95);
			MULT_96(77)<=signed(DIN_96_7)*signed(FMAP_78_96);
			MULT_97(77)<=signed(DIN_97_7)*signed(FMAP_78_97);
			MULT_98(77)<=signed(DIN_98_7)*signed(FMAP_78_98);
			MULT_99(77)<=signed(DIN_99_7)*signed(FMAP_78_99);
			MULT_100(77)<=signed(DIN_100_7)*signed(FMAP_78_100);
			MULT_101(77)<=signed(DIN_101_7)*signed(FMAP_78_101);
			MULT_102(77)<=signed(DIN_102_7)*signed(FMAP_78_102);
			MULT_103(77)<=signed(DIN_103_7)*signed(FMAP_78_103);
			MULT_104(77)<=signed(DIN_104_7)*signed(FMAP_78_104);
			MULT_105(77)<=signed(DIN_105_7)*signed(FMAP_78_105);
			MULT_106(77)<=signed(DIN_106_7)*signed(FMAP_78_106);
			MULT_107(77)<=signed(DIN_107_7)*signed(FMAP_78_107);
			MULT_108(77)<=signed(DIN_108_7)*signed(FMAP_78_108);
			MULT_109(77)<=signed(DIN_109_7)*signed(FMAP_78_109);
			MULT_110(77)<=signed(DIN_110_7)*signed(FMAP_78_110);
			MULT_111(77)<=signed(DIN_111_7)*signed(FMAP_78_111);
			MULT_112(77)<=signed(DIN_112_7)*signed(FMAP_78_112);
			MULT_113(77)<=signed(DIN_113_7)*signed(FMAP_78_113);
			MULT_114(77)<=signed(DIN_114_7)*signed(FMAP_78_114);
			MULT_115(77)<=signed(DIN_115_7)*signed(FMAP_78_115);
			MULT_116(77)<=signed(DIN_116_7)*signed(FMAP_78_116);
			MULT_117(77)<=signed(DIN_117_7)*signed(FMAP_78_117);
			MULT_118(77)<=signed(DIN_118_7)*signed(FMAP_78_118);
			MULT_119(77)<=signed(DIN_119_7)*signed(FMAP_78_119);
			MULT_120(77)<=signed(DIN_120_7)*signed(FMAP_78_120);

			MULT_1(78)<=signed(DIN_1_7)*signed(FMAP_79_1);
			MULT_2(78)<=signed(DIN_2_7)*signed(FMAP_79_2);
			MULT_3(78)<=signed(DIN_3_7)*signed(FMAP_79_3);
			MULT_4(78)<=signed(DIN_4_7)*signed(FMAP_79_4);
			MULT_5(78)<=signed(DIN_5_7)*signed(FMAP_79_5);
			MULT_6(78)<=signed(DIN_6_7)*signed(FMAP_79_6);
			MULT_7(78)<=signed(DIN_7_7)*signed(FMAP_79_7);
			MULT_8(78)<=signed(DIN_8_7)*signed(FMAP_79_8);
			MULT_9(78)<=signed(DIN_9_7)*signed(FMAP_79_9);
			MULT_10(78)<=signed(DIN_10_7)*signed(FMAP_79_10);
			MULT_11(78)<=signed(DIN_11_7)*signed(FMAP_79_11);
			MULT_12(78)<=signed(DIN_12_7)*signed(FMAP_79_12);
			MULT_13(78)<=signed(DIN_13_7)*signed(FMAP_79_13);
			MULT_14(78)<=signed(DIN_14_7)*signed(FMAP_79_14);
			MULT_15(78)<=signed(DIN_15_7)*signed(FMAP_79_15);
			MULT_16(78)<=signed(DIN_16_7)*signed(FMAP_79_16);
			MULT_17(78)<=signed(DIN_17_7)*signed(FMAP_79_17);
			MULT_18(78)<=signed(DIN_18_7)*signed(FMAP_79_18);
			MULT_19(78)<=signed(DIN_19_7)*signed(FMAP_79_19);
			MULT_20(78)<=signed(DIN_20_7)*signed(FMAP_79_20);
			MULT_21(78)<=signed(DIN_21_7)*signed(FMAP_79_21);
			MULT_22(78)<=signed(DIN_22_7)*signed(FMAP_79_22);
			MULT_23(78)<=signed(DIN_23_7)*signed(FMAP_79_23);
			MULT_24(78)<=signed(DIN_24_7)*signed(FMAP_79_24);
			MULT_25(78)<=signed(DIN_25_7)*signed(FMAP_79_25);
			MULT_26(78)<=signed(DIN_26_7)*signed(FMAP_79_26);
			MULT_27(78)<=signed(DIN_27_7)*signed(FMAP_79_27);
			MULT_28(78)<=signed(DIN_28_7)*signed(FMAP_79_28);
			MULT_29(78)<=signed(DIN_29_7)*signed(FMAP_79_29);
			MULT_30(78)<=signed(DIN_30_7)*signed(FMAP_79_30);
			MULT_31(78)<=signed(DIN_31_7)*signed(FMAP_79_31);
			MULT_32(78)<=signed(DIN_32_7)*signed(FMAP_79_32);
			MULT_33(78)<=signed(DIN_33_7)*signed(FMAP_79_33);
			MULT_34(78)<=signed(DIN_34_7)*signed(FMAP_79_34);
			MULT_35(78)<=signed(DIN_35_7)*signed(FMAP_79_35);
			MULT_36(78)<=signed(DIN_36_7)*signed(FMAP_79_36);
			MULT_37(78)<=signed(DIN_37_7)*signed(FMAP_79_37);
			MULT_38(78)<=signed(DIN_38_7)*signed(FMAP_79_38);
			MULT_39(78)<=signed(DIN_39_7)*signed(FMAP_79_39);
			MULT_40(78)<=signed(DIN_40_7)*signed(FMAP_79_40);
			MULT_41(78)<=signed(DIN_41_7)*signed(FMAP_79_41);
			MULT_42(78)<=signed(DIN_42_7)*signed(FMAP_79_42);
			MULT_43(78)<=signed(DIN_43_7)*signed(FMAP_79_43);
			MULT_44(78)<=signed(DIN_44_7)*signed(FMAP_79_44);
			MULT_45(78)<=signed(DIN_45_7)*signed(FMAP_79_45);
			MULT_46(78)<=signed(DIN_46_7)*signed(FMAP_79_46);
			MULT_47(78)<=signed(DIN_47_7)*signed(FMAP_79_47);
			MULT_48(78)<=signed(DIN_48_7)*signed(FMAP_79_48);
			MULT_49(78)<=signed(DIN_49_7)*signed(FMAP_79_49);
			MULT_50(78)<=signed(DIN_50_7)*signed(FMAP_79_50);
			MULT_51(78)<=signed(DIN_51_7)*signed(FMAP_79_51);
			MULT_52(78)<=signed(DIN_52_7)*signed(FMAP_79_52);
			MULT_53(78)<=signed(DIN_53_7)*signed(FMAP_79_53);
			MULT_54(78)<=signed(DIN_54_7)*signed(FMAP_79_54);
			MULT_55(78)<=signed(DIN_55_7)*signed(FMAP_79_55);
			MULT_56(78)<=signed(DIN_56_7)*signed(FMAP_79_56);
			MULT_57(78)<=signed(DIN_57_7)*signed(FMAP_79_57);
			MULT_58(78)<=signed(DIN_58_7)*signed(FMAP_79_58);
			MULT_59(78)<=signed(DIN_59_7)*signed(FMAP_79_59);
			MULT_60(78)<=signed(DIN_60_7)*signed(FMAP_79_60);
			MULT_61(78)<=signed(DIN_61_7)*signed(FMAP_79_61);
			MULT_62(78)<=signed(DIN_62_7)*signed(FMAP_79_62);
			MULT_63(78)<=signed(DIN_63_7)*signed(FMAP_79_63);
			MULT_64(78)<=signed(DIN_64_7)*signed(FMAP_79_64);
			MULT_65(78)<=signed(DIN_65_7)*signed(FMAP_79_65);
			MULT_66(78)<=signed(DIN_66_7)*signed(FMAP_79_66);
			MULT_67(78)<=signed(DIN_67_7)*signed(FMAP_79_67);
			MULT_68(78)<=signed(DIN_68_7)*signed(FMAP_79_68);
			MULT_69(78)<=signed(DIN_69_7)*signed(FMAP_79_69);
			MULT_70(78)<=signed(DIN_70_7)*signed(FMAP_79_70);
			MULT_71(78)<=signed(DIN_71_7)*signed(FMAP_79_71);
			MULT_72(78)<=signed(DIN_72_7)*signed(FMAP_79_72);
			MULT_73(78)<=signed(DIN_73_7)*signed(FMAP_79_73);
			MULT_74(78)<=signed(DIN_74_7)*signed(FMAP_79_74);
			MULT_75(78)<=signed(DIN_75_7)*signed(FMAP_79_75);
			MULT_76(78)<=signed(DIN_76_7)*signed(FMAP_79_76);
			MULT_77(78)<=signed(DIN_77_7)*signed(FMAP_79_77);
			MULT_78(78)<=signed(DIN_78_7)*signed(FMAP_79_78);
			MULT_79(78)<=signed(DIN_79_7)*signed(FMAP_79_79);
			MULT_80(78)<=signed(DIN_80_7)*signed(FMAP_79_80);
			MULT_81(78)<=signed(DIN_81_7)*signed(FMAP_79_81);
			MULT_82(78)<=signed(DIN_82_7)*signed(FMAP_79_82);
			MULT_83(78)<=signed(DIN_83_7)*signed(FMAP_79_83);
			MULT_84(78)<=signed(DIN_84_7)*signed(FMAP_79_84);
			MULT_85(78)<=signed(DIN_85_7)*signed(FMAP_79_85);
			MULT_86(78)<=signed(DIN_86_7)*signed(FMAP_79_86);
			MULT_87(78)<=signed(DIN_87_7)*signed(FMAP_79_87);
			MULT_88(78)<=signed(DIN_88_7)*signed(FMAP_79_88);
			MULT_89(78)<=signed(DIN_89_7)*signed(FMAP_79_89);
			MULT_90(78)<=signed(DIN_90_7)*signed(FMAP_79_90);
			MULT_91(78)<=signed(DIN_91_7)*signed(FMAP_79_91);
			MULT_92(78)<=signed(DIN_92_7)*signed(FMAP_79_92);
			MULT_93(78)<=signed(DIN_93_7)*signed(FMAP_79_93);
			MULT_94(78)<=signed(DIN_94_7)*signed(FMAP_79_94);
			MULT_95(78)<=signed(DIN_95_7)*signed(FMAP_79_95);
			MULT_96(78)<=signed(DIN_96_7)*signed(FMAP_79_96);
			MULT_97(78)<=signed(DIN_97_7)*signed(FMAP_79_97);
			MULT_98(78)<=signed(DIN_98_7)*signed(FMAP_79_98);
			MULT_99(78)<=signed(DIN_99_7)*signed(FMAP_79_99);
			MULT_100(78)<=signed(DIN_100_7)*signed(FMAP_79_100);
			MULT_101(78)<=signed(DIN_101_7)*signed(FMAP_79_101);
			MULT_102(78)<=signed(DIN_102_7)*signed(FMAP_79_102);
			MULT_103(78)<=signed(DIN_103_7)*signed(FMAP_79_103);
			MULT_104(78)<=signed(DIN_104_7)*signed(FMAP_79_104);
			MULT_105(78)<=signed(DIN_105_7)*signed(FMAP_79_105);
			MULT_106(78)<=signed(DIN_106_7)*signed(FMAP_79_106);
			MULT_107(78)<=signed(DIN_107_7)*signed(FMAP_79_107);
			MULT_108(78)<=signed(DIN_108_7)*signed(FMAP_79_108);
			MULT_109(78)<=signed(DIN_109_7)*signed(FMAP_79_109);
			MULT_110(78)<=signed(DIN_110_7)*signed(FMAP_79_110);
			MULT_111(78)<=signed(DIN_111_7)*signed(FMAP_79_111);
			MULT_112(78)<=signed(DIN_112_7)*signed(FMAP_79_112);
			MULT_113(78)<=signed(DIN_113_7)*signed(FMAP_79_113);
			MULT_114(78)<=signed(DIN_114_7)*signed(FMAP_79_114);
			MULT_115(78)<=signed(DIN_115_7)*signed(FMAP_79_115);
			MULT_116(78)<=signed(DIN_116_7)*signed(FMAP_79_116);
			MULT_117(78)<=signed(DIN_117_7)*signed(FMAP_79_117);
			MULT_118(78)<=signed(DIN_118_7)*signed(FMAP_79_118);
			MULT_119(78)<=signed(DIN_119_7)*signed(FMAP_79_119);
			MULT_120(78)<=signed(DIN_120_7)*signed(FMAP_79_120);

			MULT_1(79)<=signed(DIN_1_7)*signed(FMAP_80_1);
			MULT_2(79)<=signed(DIN_2_7)*signed(FMAP_80_2);
			MULT_3(79)<=signed(DIN_3_7)*signed(FMAP_80_3);
			MULT_4(79)<=signed(DIN_4_7)*signed(FMAP_80_4);
			MULT_5(79)<=signed(DIN_5_7)*signed(FMAP_80_5);
			MULT_6(79)<=signed(DIN_6_7)*signed(FMAP_80_6);
			MULT_7(79)<=signed(DIN_7_7)*signed(FMAP_80_7);
			MULT_8(79)<=signed(DIN_8_7)*signed(FMAP_80_8);
			MULT_9(79)<=signed(DIN_9_7)*signed(FMAP_80_9);
			MULT_10(79)<=signed(DIN_10_7)*signed(FMAP_80_10);
			MULT_11(79)<=signed(DIN_11_7)*signed(FMAP_80_11);
			MULT_12(79)<=signed(DIN_12_7)*signed(FMAP_80_12);
			MULT_13(79)<=signed(DIN_13_7)*signed(FMAP_80_13);
			MULT_14(79)<=signed(DIN_14_7)*signed(FMAP_80_14);
			MULT_15(79)<=signed(DIN_15_7)*signed(FMAP_80_15);
			MULT_16(79)<=signed(DIN_16_7)*signed(FMAP_80_16);
			MULT_17(79)<=signed(DIN_17_7)*signed(FMAP_80_17);
			MULT_18(79)<=signed(DIN_18_7)*signed(FMAP_80_18);
			MULT_19(79)<=signed(DIN_19_7)*signed(FMAP_80_19);
			MULT_20(79)<=signed(DIN_20_7)*signed(FMAP_80_20);
			MULT_21(79)<=signed(DIN_21_7)*signed(FMAP_80_21);
			MULT_22(79)<=signed(DIN_22_7)*signed(FMAP_80_22);
			MULT_23(79)<=signed(DIN_23_7)*signed(FMAP_80_23);
			MULT_24(79)<=signed(DIN_24_7)*signed(FMAP_80_24);
			MULT_25(79)<=signed(DIN_25_7)*signed(FMAP_80_25);
			MULT_26(79)<=signed(DIN_26_7)*signed(FMAP_80_26);
			MULT_27(79)<=signed(DIN_27_7)*signed(FMAP_80_27);
			MULT_28(79)<=signed(DIN_28_7)*signed(FMAP_80_28);
			MULT_29(79)<=signed(DIN_29_7)*signed(FMAP_80_29);
			MULT_30(79)<=signed(DIN_30_7)*signed(FMAP_80_30);
			MULT_31(79)<=signed(DIN_31_7)*signed(FMAP_80_31);
			MULT_32(79)<=signed(DIN_32_7)*signed(FMAP_80_32);
			MULT_33(79)<=signed(DIN_33_7)*signed(FMAP_80_33);
			MULT_34(79)<=signed(DIN_34_7)*signed(FMAP_80_34);
			MULT_35(79)<=signed(DIN_35_7)*signed(FMAP_80_35);
			MULT_36(79)<=signed(DIN_36_7)*signed(FMAP_80_36);
			MULT_37(79)<=signed(DIN_37_7)*signed(FMAP_80_37);
			MULT_38(79)<=signed(DIN_38_7)*signed(FMAP_80_38);
			MULT_39(79)<=signed(DIN_39_7)*signed(FMAP_80_39);
			MULT_40(79)<=signed(DIN_40_7)*signed(FMAP_80_40);
			MULT_41(79)<=signed(DIN_41_7)*signed(FMAP_80_41);
			MULT_42(79)<=signed(DIN_42_7)*signed(FMAP_80_42);
			MULT_43(79)<=signed(DIN_43_7)*signed(FMAP_80_43);
			MULT_44(79)<=signed(DIN_44_7)*signed(FMAP_80_44);
			MULT_45(79)<=signed(DIN_45_7)*signed(FMAP_80_45);
			MULT_46(79)<=signed(DIN_46_7)*signed(FMAP_80_46);
			MULT_47(79)<=signed(DIN_47_7)*signed(FMAP_80_47);
			MULT_48(79)<=signed(DIN_48_7)*signed(FMAP_80_48);
			MULT_49(79)<=signed(DIN_49_7)*signed(FMAP_80_49);
			MULT_50(79)<=signed(DIN_50_7)*signed(FMAP_80_50);
			MULT_51(79)<=signed(DIN_51_7)*signed(FMAP_80_51);
			MULT_52(79)<=signed(DIN_52_7)*signed(FMAP_80_52);
			MULT_53(79)<=signed(DIN_53_7)*signed(FMAP_80_53);
			MULT_54(79)<=signed(DIN_54_7)*signed(FMAP_80_54);
			MULT_55(79)<=signed(DIN_55_7)*signed(FMAP_80_55);
			MULT_56(79)<=signed(DIN_56_7)*signed(FMAP_80_56);
			MULT_57(79)<=signed(DIN_57_7)*signed(FMAP_80_57);
			MULT_58(79)<=signed(DIN_58_7)*signed(FMAP_80_58);
			MULT_59(79)<=signed(DIN_59_7)*signed(FMAP_80_59);
			MULT_60(79)<=signed(DIN_60_7)*signed(FMAP_80_60);
			MULT_61(79)<=signed(DIN_61_7)*signed(FMAP_80_61);
			MULT_62(79)<=signed(DIN_62_7)*signed(FMAP_80_62);
			MULT_63(79)<=signed(DIN_63_7)*signed(FMAP_80_63);
			MULT_64(79)<=signed(DIN_64_7)*signed(FMAP_80_64);
			MULT_65(79)<=signed(DIN_65_7)*signed(FMAP_80_65);
			MULT_66(79)<=signed(DIN_66_7)*signed(FMAP_80_66);
			MULT_67(79)<=signed(DIN_67_7)*signed(FMAP_80_67);
			MULT_68(79)<=signed(DIN_68_7)*signed(FMAP_80_68);
			MULT_69(79)<=signed(DIN_69_7)*signed(FMAP_80_69);
			MULT_70(79)<=signed(DIN_70_7)*signed(FMAP_80_70);
			MULT_71(79)<=signed(DIN_71_7)*signed(FMAP_80_71);
			MULT_72(79)<=signed(DIN_72_7)*signed(FMAP_80_72);
			MULT_73(79)<=signed(DIN_73_7)*signed(FMAP_80_73);
			MULT_74(79)<=signed(DIN_74_7)*signed(FMAP_80_74);
			MULT_75(79)<=signed(DIN_75_7)*signed(FMAP_80_75);
			MULT_76(79)<=signed(DIN_76_7)*signed(FMAP_80_76);
			MULT_77(79)<=signed(DIN_77_7)*signed(FMAP_80_77);
			MULT_78(79)<=signed(DIN_78_7)*signed(FMAP_80_78);
			MULT_79(79)<=signed(DIN_79_7)*signed(FMAP_80_79);
			MULT_80(79)<=signed(DIN_80_7)*signed(FMAP_80_80);
			MULT_81(79)<=signed(DIN_81_7)*signed(FMAP_80_81);
			MULT_82(79)<=signed(DIN_82_7)*signed(FMAP_80_82);
			MULT_83(79)<=signed(DIN_83_7)*signed(FMAP_80_83);
			MULT_84(79)<=signed(DIN_84_7)*signed(FMAP_80_84);
			MULT_85(79)<=signed(DIN_85_7)*signed(FMAP_80_85);
			MULT_86(79)<=signed(DIN_86_7)*signed(FMAP_80_86);
			MULT_87(79)<=signed(DIN_87_7)*signed(FMAP_80_87);
			MULT_88(79)<=signed(DIN_88_7)*signed(FMAP_80_88);
			MULT_89(79)<=signed(DIN_89_7)*signed(FMAP_80_89);
			MULT_90(79)<=signed(DIN_90_7)*signed(FMAP_80_90);
			MULT_91(79)<=signed(DIN_91_7)*signed(FMAP_80_91);
			MULT_92(79)<=signed(DIN_92_7)*signed(FMAP_80_92);
			MULT_93(79)<=signed(DIN_93_7)*signed(FMAP_80_93);
			MULT_94(79)<=signed(DIN_94_7)*signed(FMAP_80_94);
			MULT_95(79)<=signed(DIN_95_7)*signed(FMAP_80_95);
			MULT_96(79)<=signed(DIN_96_7)*signed(FMAP_80_96);
			MULT_97(79)<=signed(DIN_97_7)*signed(FMAP_80_97);
			MULT_98(79)<=signed(DIN_98_7)*signed(FMAP_80_98);
			MULT_99(79)<=signed(DIN_99_7)*signed(FMAP_80_99);
			MULT_100(79)<=signed(DIN_100_7)*signed(FMAP_80_100);
			MULT_101(79)<=signed(DIN_101_7)*signed(FMAP_80_101);
			MULT_102(79)<=signed(DIN_102_7)*signed(FMAP_80_102);
			MULT_103(79)<=signed(DIN_103_7)*signed(FMAP_80_103);
			MULT_104(79)<=signed(DIN_104_7)*signed(FMAP_80_104);
			MULT_105(79)<=signed(DIN_105_7)*signed(FMAP_80_105);
			MULT_106(79)<=signed(DIN_106_7)*signed(FMAP_80_106);
			MULT_107(79)<=signed(DIN_107_7)*signed(FMAP_80_107);
			MULT_108(79)<=signed(DIN_108_7)*signed(FMAP_80_108);
			MULT_109(79)<=signed(DIN_109_7)*signed(FMAP_80_109);
			MULT_110(79)<=signed(DIN_110_7)*signed(FMAP_80_110);
			MULT_111(79)<=signed(DIN_111_7)*signed(FMAP_80_111);
			MULT_112(79)<=signed(DIN_112_7)*signed(FMAP_80_112);
			MULT_113(79)<=signed(DIN_113_7)*signed(FMAP_80_113);
			MULT_114(79)<=signed(DIN_114_7)*signed(FMAP_80_114);
			MULT_115(79)<=signed(DIN_115_7)*signed(FMAP_80_115);
			MULT_116(79)<=signed(DIN_116_7)*signed(FMAP_80_116);
			MULT_117(79)<=signed(DIN_117_7)*signed(FMAP_80_117);
			MULT_118(79)<=signed(DIN_118_7)*signed(FMAP_80_118);
			MULT_119(79)<=signed(DIN_119_7)*signed(FMAP_80_119);
			MULT_120(79)<=signed(DIN_120_7)*signed(FMAP_80_120);

			MULT_1(80)<=signed(DIN_1_7)*signed(FMAP_81_1);
			MULT_2(80)<=signed(DIN_2_7)*signed(FMAP_81_2);
			MULT_3(80)<=signed(DIN_3_7)*signed(FMAP_81_3);
			MULT_4(80)<=signed(DIN_4_7)*signed(FMAP_81_4);
			MULT_5(80)<=signed(DIN_5_7)*signed(FMAP_81_5);
			MULT_6(80)<=signed(DIN_6_7)*signed(FMAP_81_6);
			MULT_7(80)<=signed(DIN_7_7)*signed(FMAP_81_7);
			MULT_8(80)<=signed(DIN_8_7)*signed(FMAP_81_8);
			MULT_9(80)<=signed(DIN_9_7)*signed(FMAP_81_9);
			MULT_10(80)<=signed(DIN_10_7)*signed(FMAP_81_10);
			MULT_11(80)<=signed(DIN_11_7)*signed(FMAP_81_11);
			MULT_12(80)<=signed(DIN_12_7)*signed(FMAP_81_12);
			MULT_13(80)<=signed(DIN_13_7)*signed(FMAP_81_13);
			MULT_14(80)<=signed(DIN_14_7)*signed(FMAP_81_14);
			MULT_15(80)<=signed(DIN_15_7)*signed(FMAP_81_15);
			MULT_16(80)<=signed(DIN_16_7)*signed(FMAP_81_16);
			MULT_17(80)<=signed(DIN_17_7)*signed(FMAP_81_17);
			MULT_18(80)<=signed(DIN_18_7)*signed(FMAP_81_18);
			MULT_19(80)<=signed(DIN_19_7)*signed(FMAP_81_19);
			MULT_20(80)<=signed(DIN_20_7)*signed(FMAP_81_20);
			MULT_21(80)<=signed(DIN_21_7)*signed(FMAP_81_21);
			MULT_22(80)<=signed(DIN_22_7)*signed(FMAP_81_22);
			MULT_23(80)<=signed(DIN_23_7)*signed(FMAP_81_23);
			MULT_24(80)<=signed(DIN_24_7)*signed(FMAP_81_24);
			MULT_25(80)<=signed(DIN_25_7)*signed(FMAP_81_25);
			MULT_26(80)<=signed(DIN_26_7)*signed(FMAP_81_26);
			MULT_27(80)<=signed(DIN_27_7)*signed(FMAP_81_27);
			MULT_28(80)<=signed(DIN_28_7)*signed(FMAP_81_28);
			MULT_29(80)<=signed(DIN_29_7)*signed(FMAP_81_29);
			MULT_30(80)<=signed(DIN_30_7)*signed(FMAP_81_30);
			MULT_31(80)<=signed(DIN_31_7)*signed(FMAP_81_31);
			MULT_32(80)<=signed(DIN_32_7)*signed(FMAP_81_32);
			MULT_33(80)<=signed(DIN_33_7)*signed(FMAP_81_33);
			MULT_34(80)<=signed(DIN_34_7)*signed(FMAP_81_34);
			MULT_35(80)<=signed(DIN_35_7)*signed(FMAP_81_35);
			MULT_36(80)<=signed(DIN_36_7)*signed(FMAP_81_36);
			MULT_37(80)<=signed(DIN_37_7)*signed(FMAP_81_37);
			MULT_38(80)<=signed(DIN_38_7)*signed(FMAP_81_38);
			MULT_39(80)<=signed(DIN_39_7)*signed(FMAP_81_39);
			MULT_40(80)<=signed(DIN_40_7)*signed(FMAP_81_40);
			MULT_41(80)<=signed(DIN_41_7)*signed(FMAP_81_41);
			MULT_42(80)<=signed(DIN_42_7)*signed(FMAP_81_42);
			MULT_43(80)<=signed(DIN_43_7)*signed(FMAP_81_43);
			MULT_44(80)<=signed(DIN_44_7)*signed(FMAP_81_44);
			MULT_45(80)<=signed(DIN_45_7)*signed(FMAP_81_45);
			MULT_46(80)<=signed(DIN_46_7)*signed(FMAP_81_46);
			MULT_47(80)<=signed(DIN_47_7)*signed(FMAP_81_47);
			MULT_48(80)<=signed(DIN_48_7)*signed(FMAP_81_48);
			MULT_49(80)<=signed(DIN_49_7)*signed(FMAP_81_49);
			MULT_50(80)<=signed(DIN_50_7)*signed(FMAP_81_50);
			MULT_51(80)<=signed(DIN_51_7)*signed(FMAP_81_51);
			MULT_52(80)<=signed(DIN_52_7)*signed(FMAP_81_52);
			MULT_53(80)<=signed(DIN_53_7)*signed(FMAP_81_53);
			MULT_54(80)<=signed(DIN_54_7)*signed(FMAP_81_54);
			MULT_55(80)<=signed(DIN_55_7)*signed(FMAP_81_55);
			MULT_56(80)<=signed(DIN_56_7)*signed(FMAP_81_56);
			MULT_57(80)<=signed(DIN_57_7)*signed(FMAP_81_57);
			MULT_58(80)<=signed(DIN_58_7)*signed(FMAP_81_58);
			MULT_59(80)<=signed(DIN_59_7)*signed(FMAP_81_59);
			MULT_60(80)<=signed(DIN_60_7)*signed(FMAP_81_60);
			MULT_61(80)<=signed(DIN_61_7)*signed(FMAP_81_61);
			MULT_62(80)<=signed(DIN_62_7)*signed(FMAP_81_62);
			MULT_63(80)<=signed(DIN_63_7)*signed(FMAP_81_63);
			MULT_64(80)<=signed(DIN_64_7)*signed(FMAP_81_64);
			MULT_65(80)<=signed(DIN_65_7)*signed(FMAP_81_65);
			MULT_66(80)<=signed(DIN_66_7)*signed(FMAP_81_66);
			MULT_67(80)<=signed(DIN_67_7)*signed(FMAP_81_67);
			MULT_68(80)<=signed(DIN_68_7)*signed(FMAP_81_68);
			MULT_69(80)<=signed(DIN_69_7)*signed(FMAP_81_69);
			MULT_70(80)<=signed(DIN_70_7)*signed(FMAP_81_70);
			MULT_71(80)<=signed(DIN_71_7)*signed(FMAP_81_71);
			MULT_72(80)<=signed(DIN_72_7)*signed(FMAP_81_72);
			MULT_73(80)<=signed(DIN_73_7)*signed(FMAP_81_73);
			MULT_74(80)<=signed(DIN_74_7)*signed(FMAP_81_74);
			MULT_75(80)<=signed(DIN_75_7)*signed(FMAP_81_75);
			MULT_76(80)<=signed(DIN_76_7)*signed(FMAP_81_76);
			MULT_77(80)<=signed(DIN_77_7)*signed(FMAP_81_77);
			MULT_78(80)<=signed(DIN_78_7)*signed(FMAP_81_78);
			MULT_79(80)<=signed(DIN_79_7)*signed(FMAP_81_79);
			MULT_80(80)<=signed(DIN_80_7)*signed(FMAP_81_80);
			MULT_81(80)<=signed(DIN_81_7)*signed(FMAP_81_81);
			MULT_82(80)<=signed(DIN_82_7)*signed(FMAP_81_82);
			MULT_83(80)<=signed(DIN_83_7)*signed(FMAP_81_83);
			MULT_84(80)<=signed(DIN_84_7)*signed(FMAP_81_84);
			MULT_85(80)<=signed(DIN_85_7)*signed(FMAP_81_85);
			MULT_86(80)<=signed(DIN_86_7)*signed(FMAP_81_86);
			MULT_87(80)<=signed(DIN_87_7)*signed(FMAP_81_87);
			MULT_88(80)<=signed(DIN_88_7)*signed(FMAP_81_88);
			MULT_89(80)<=signed(DIN_89_7)*signed(FMAP_81_89);
			MULT_90(80)<=signed(DIN_90_7)*signed(FMAP_81_90);
			MULT_91(80)<=signed(DIN_91_7)*signed(FMAP_81_91);
			MULT_92(80)<=signed(DIN_92_7)*signed(FMAP_81_92);
			MULT_93(80)<=signed(DIN_93_7)*signed(FMAP_81_93);
			MULT_94(80)<=signed(DIN_94_7)*signed(FMAP_81_94);
			MULT_95(80)<=signed(DIN_95_7)*signed(FMAP_81_95);
			MULT_96(80)<=signed(DIN_96_7)*signed(FMAP_81_96);
			MULT_97(80)<=signed(DIN_97_7)*signed(FMAP_81_97);
			MULT_98(80)<=signed(DIN_98_7)*signed(FMAP_81_98);
			MULT_99(80)<=signed(DIN_99_7)*signed(FMAP_81_99);
			MULT_100(80)<=signed(DIN_100_7)*signed(FMAP_81_100);
			MULT_101(80)<=signed(DIN_101_7)*signed(FMAP_81_101);
			MULT_102(80)<=signed(DIN_102_7)*signed(FMAP_81_102);
			MULT_103(80)<=signed(DIN_103_7)*signed(FMAP_81_103);
			MULT_104(80)<=signed(DIN_104_7)*signed(FMAP_81_104);
			MULT_105(80)<=signed(DIN_105_7)*signed(FMAP_81_105);
			MULT_106(80)<=signed(DIN_106_7)*signed(FMAP_81_106);
			MULT_107(80)<=signed(DIN_107_7)*signed(FMAP_81_107);
			MULT_108(80)<=signed(DIN_108_7)*signed(FMAP_81_108);
			MULT_109(80)<=signed(DIN_109_7)*signed(FMAP_81_109);
			MULT_110(80)<=signed(DIN_110_7)*signed(FMAP_81_110);
			MULT_111(80)<=signed(DIN_111_7)*signed(FMAP_81_111);
			MULT_112(80)<=signed(DIN_112_7)*signed(FMAP_81_112);
			MULT_113(80)<=signed(DIN_113_7)*signed(FMAP_81_113);
			MULT_114(80)<=signed(DIN_114_7)*signed(FMAP_81_114);
			MULT_115(80)<=signed(DIN_115_7)*signed(FMAP_81_115);
			MULT_116(80)<=signed(DIN_116_7)*signed(FMAP_81_116);
			MULT_117(80)<=signed(DIN_117_7)*signed(FMAP_81_117);
			MULT_118(80)<=signed(DIN_118_7)*signed(FMAP_81_118);
			MULT_119(80)<=signed(DIN_119_7)*signed(FMAP_81_119);
			MULT_120(80)<=signed(DIN_120_7)*signed(FMAP_81_120);

			MULT_1(81)<=signed(DIN_1_7)*signed(FMAP_82_1);
			MULT_2(81)<=signed(DIN_2_7)*signed(FMAP_82_2);
			MULT_3(81)<=signed(DIN_3_7)*signed(FMAP_82_3);
			MULT_4(81)<=signed(DIN_4_7)*signed(FMAP_82_4);
			MULT_5(81)<=signed(DIN_5_7)*signed(FMAP_82_5);
			MULT_6(81)<=signed(DIN_6_7)*signed(FMAP_82_6);
			MULT_7(81)<=signed(DIN_7_7)*signed(FMAP_82_7);
			MULT_8(81)<=signed(DIN_8_7)*signed(FMAP_82_8);
			MULT_9(81)<=signed(DIN_9_7)*signed(FMAP_82_9);
			MULT_10(81)<=signed(DIN_10_7)*signed(FMAP_82_10);
			MULT_11(81)<=signed(DIN_11_7)*signed(FMAP_82_11);
			MULT_12(81)<=signed(DIN_12_7)*signed(FMAP_82_12);
			MULT_13(81)<=signed(DIN_13_7)*signed(FMAP_82_13);
			MULT_14(81)<=signed(DIN_14_7)*signed(FMAP_82_14);
			MULT_15(81)<=signed(DIN_15_7)*signed(FMAP_82_15);
			MULT_16(81)<=signed(DIN_16_7)*signed(FMAP_82_16);
			MULT_17(81)<=signed(DIN_17_7)*signed(FMAP_82_17);
			MULT_18(81)<=signed(DIN_18_7)*signed(FMAP_82_18);
			MULT_19(81)<=signed(DIN_19_7)*signed(FMAP_82_19);
			MULT_20(81)<=signed(DIN_20_7)*signed(FMAP_82_20);
			MULT_21(81)<=signed(DIN_21_7)*signed(FMAP_82_21);
			MULT_22(81)<=signed(DIN_22_7)*signed(FMAP_82_22);
			MULT_23(81)<=signed(DIN_23_7)*signed(FMAP_82_23);
			MULT_24(81)<=signed(DIN_24_7)*signed(FMAP_82_24);
			MULT_25(81)<=signed(DIN_25_7)*signed(FMAP_82_25);
			MULT_26(81)<=signed(DIN_26_7)*signed(FMAP_82_26);
			MULT_27(81)<=signed(DIN_27_7)*signed(FMAP_82_27);
			MULT_28(81)<=signed(DIN_28_7)*signed(FMAP_82_28);
			MULT_29(81)<=signed(DIN_29_7)*signed(FMAP_82_29);
			MULT_30(81)<=signed(DIN_30_7)*signed(FMAP_82_30);
			MULT_31(81)<=signed(DIN_31_7)*signed(FMAP_82_31);
			MULT_32(81)<=signed(DIN_32_7)*signed(FMAP_82_32);
			MULT_33(81)<=signed(DIN_33_7)*signed(FMAP_82_33);
			MULT_34(81)<=signed(DIN_34_7)*signed(FMAP_82_34);
			MULT_35(81)<=signed(DIN_35_7)*signed(FMAP_82_35);
			MULT_36(81)<=signed(DIN_36_7)*signed(FMAP_82_36);
			MULT_37(81)<=signed(DIN_37_7)*signed(FMAP_82_37);
			MULT_38(81)<=signed(DIN_38_7)*signed(FMAP_82_38);
			MULT_39(81)<=signed(DIN_39_7)*signed(FMAP_82_39);
			MULT_40(81)<=signed(DIN_40_7)*signed(FMAP_82_40);
			MULT_41(81)<=signed(DIN_41_7)*signed(FMAP_82_41);
			MULT_42(81)<=signed(DIN_42_7)*signed(FMAP_82_42);
			MULT_43(81)<=signed(DIN_43_7)*signed(FMAP_82_43);
			MULT_44(81)<=signed(DIN_44_7)*signed(FMAP_82_44);
			MULT_45(81)<=signed(DIN_45_7)*signed(FMAP_82_45);
			MULT_46(81)<=signed(DIN_46_7)*signed(FMAP_82_46);
			MULT_47(81)<=signed(DIN_47_7)*signed(FMAP_82_47);
			MULT_48(81)<=signed(DIN_48_7)*signed(FMAP_82_48);
			MULT_49(81)<=signed(DIN_49_7)*signed(FMAP_82_49);
			MULT_50(81)<=signed(DIN_50_7)*signed(FMAP_82_50);
			MULT_51(81)<=signed(DIN_51_7)*signed(FMAP_82_51);
			MULT_52(81)<=signed(DIN_52_7)*signed(FMAP_82_52);
			MULT_53(81)<=signed(DIN_53_7)*signed(FMAP_82_53);
			MULT_54(81)<=signed(DIN_54_7)*signed(FMAP_82_54);
			MULT_55(81)<=signed(DIN_55_7)*signed(FMAP_82_55);
			MULT_56(81)<=signed(DIN_56_7)*signed(FMAP_82_56);
			MULT_57(81)<=signed(DIN_57_7)*signed(FMAP_82_57);
			MULT_58(81)<=signed(DIN_58_7)*signed(FMAP_82_58);
			MULT_59(81)<=signed(DIN_59_7)*signed(FMAP_82_59);
			MULT_60(81)<=signed(DIN_60_7)*signed(FMAP_82_60);
			MULT_61(81)<=signed(DIN_61_7)*signed(FMAP_82_61);
			MULT_62(81)<=signed(DIN_62_7)*signed(FMAP_82_62);
			MULT_63(81)<=signed(DIN_63_7)*signed(FMAP_82_63);
			MULT_64(81)<=signed(DIN_64_7)*signed(FMAP_82_64);
			MULT_65(81)<=signed(DIN_65_7)*signed(FMAP_82_65);
			MULT_66(81)<=signed(DIN_66_7)*signed(FMAP_82_66);
			MULT_67(81)<=signed(DIN_67_7)*signed(FMAP_82_67);
			MULT_68(81)<=signed(DIN_68_7)*signed(FMAP_82_68);
			MULT_69(81)<=signed(DIN_69_7)*signed(FMAP_82_69);
			MULT_70(81)<=signed(DIN_70_7)*signed(FMAP_82_70);
			MULT_71(81)<=signed(DIN_71_7)*signed(FMAP_82_71);
			MULT_72(81)<=signed(DIN_72_7)*signed(FMAP_82_72);
			MULT_73(81)<=signed(DIN_73_7)*signed(FMAP_82_73);
			MULT_74(81)<=signed(DIN_74_7)*signed(FMAP_82_74);
			MULT_75(81)<=signed(DIN_75_7)*signed(FMAP_82_75);
			MULT_76(81)<=signed(DIN_76_7)*signed(FMAP_82_76);
			MULT_77(81)<=signed(DIN_77_7)*signed(FMAP_82_77);
			MULT_78(81)<=signed(DIN_78_7)*signed(FMAP_82_78);
			MULT_79(81)<=signed(DIN_79_7)*signed(FMAP_82_79);
			MULT_80(81)<=signed(DIN_80_7)*signed(FMAP_82_80);
			MULT_81(81)<=signed(DIN_81_7)*signed(FMAP_82_81);
			MULT_82(81)<=signed(DIN_82_7)*signed(FMAP_82_82);
			MULT_83(81)<=signed(DIN_83_7)*signed(FMAP_82_83);
			MULT_84(81)<=signed(DIN_84_7)*signed(FMAP_82_84);
			MULT_85(81)<=signed(DIN_85_7)*signed(FMAP_82_85);
			MULT_86(81)<=signed(DIN_86_7)*signed(FMAP_82_86);
			MULT_87(81)<=signed(DIN_87_7)*signed(FMAP_82_87);
			MULT_88(81)<=signed(DIN_88_7)*signed(FMAP_82_88);
			MULT_89(81)<=signed(DIN_89_7)*signed(FMAP_82_89);
			MULT_90(81)<=signed(DIN_90_7)*signed(FMAP_82_90);
			MULT_91(81)<=signed(DIN_91_7)*signed(FMAP_82_91);
			MULT_92(81)<=signed(DIN_92_7)*signed(FMAP_82_92);
			MULT_93(81)<=signed(DIN_93_7)*signed(FMAP_82_93);
			MULT_94(81)<=signed(DIN_94_7)*signed(FMAP_82_94);
			MULT_95(81)<=signed(DIN_95_7)*signed(FMAP_82_95);
			MULT_96(81)<=signed(DIN_96_7)*signed(FMAP_82_96);
			MULT_97(81)<=signed(DIN_97_7)*signed(FMAP_82_97);
			MULT_98(81)<=signed(DIN_98_7)*signed(FMAP_82_98);
			MULT_99(81)<=signed(DIN_99_7)*signed(FMAP_82_99);
			MULT_100(81)<=signed(DIN_100_7)*signed(FMAP_82_100);
			MULT_101(81)<=signed(DIN_101_7)*signed(FMAP_82_101);
			MULT_102(81)<=signed(DIN_102_7)*signed(FMAP_82_102);
			MULT_103(81)<=signed(DIN_103_7)*signed(FMAP_82_103);
			MULT_104(81)<=signed(DIN_104_7)*signed(FMAP_82_104);
			MULT_105(81)<=signed(DIN_105_7)*signed(FMAP_82_105);
			MULT_106(81)<=signed(DIN_106_7)*signed(FMAP_82_106);
			MULT_107(81)<=signed(DIN_107_7)*signed(FMAP_82_107);
			MULT_108(81)<=signed(DIN_108_7)*signed(FMAP_82_108);
			MULT_109(81)<=signed(DIN_109_7)*signed(FMAP_82_109);
			MULT_110(81)<=signed(DIN_110_7)*signed(FMAP_82_110);
			MULT_111(81)<=signed(DIN_111_7)*signed(FMAP_82_111);
			MULT_112(81)<=signed(DIN_112_7)*signed(FMAP_82_112);
			MULT_113(81)<=signed(DIN_113_7)*signed(FMAP_82_113);
			MULT_114(81)<=signed(DIN_114_7)*signed(FMAP_82_114);
			MULT_115(81)<=signed(DIN_115_7)*signed(FMAP_82_115);
			MULT_116(81)<=signed(DIN_116_7)*signed(FMAP_82_116);
			MULT_117(81)<=signed(DIN_117_7)*signed(FMAP_82_117);
			MULT_118(81)<=signed(DIN_118_7)*signed(FMAP_82_118);
			MULT_119(81)<=signed(DIN_119_7)*signed(FMAP_82_119);
			MULT_120(81)<=signed(DIN_120_7)*signed(FMAP_82_120);

			MULT_1(82)<=signed(DIN_1_7)*signed(FMAP_83_1);
			MULT_2(82)<=signed(DIN_2_7)*signed(FMAP_83_2);
			MULT_3(82)<=signed(DIN_3_7)*signed(FMAP_83_3);
			MULT_4(82)<=signed(DIN_4_7)*signed(FMAP_83_4);
			MULT_5(82)<=signed(DIN_5_7)*signed(FMAP_83_5);
			MULT_6(82)<=signed(DIN_6_7)*signed(FMAP_83_6);
			MULT_7(82)<=signed(DIN_7_7)*signed(FMAP_83_7);
			MULT_8(82)<=signed(DIN_8_7)*signed(FMAP_83_8);
			MULT_9(82)<=signed(DIN_9_7)*signed(FMAP_83_9);
			MULT_10(82)<=signed(DIN_10_7)*signed(FMAP_83_10);
			MULT_11(82)<=signed(DIN_11_7)*signed(FMAP_83_11);
			MULT_12(82)<=signed(DIN_12_7)*signed(FMAP_83_12);
			MULT_13(82)<=signed(DIN_13_7)*signed(FMAP_83_13);
			MULT_14(82)<=signed(DIN_14_7)*signed(FMAP_83_14);
			MULT_15(82)<=signed(DIN_15_7)*signed(FMAP_83_15);
			MULT_16(82)<=signed(DIN_16_7)*signed(FMAP_83_16);
			MULT_17(82)<=signed(DIN_17_7)*signed(FMAP_83_17);
			MULT_18(82)<=signed(DIN_18_7)*signed(FMAP_83_18);
			MULT_19(82)<=signed(DIN_19_7)*signed(FMAP_83_19);
			MULT_20(82)<=signed(DIN_20_7)*signed(FMAP_83_20);
			MULT_21(82)<=signed(DIN_21_7)*signed(FMAP_83_21);
			MULT_22(82)<=signed(DIN_22_7)*signed(FMAP_83_22);
			MULT_23(82)<=signed(DIN_23_7)*signed(FMAP_83_23);
			MULT_24(82)<=signed(DIN_24_7)*signed(FMAP_83_24);
			MULT_25(82)<=signed(DIN_25_7)*signed(FMAP_83_25);
			MULT_26(82)<=signed(DIN_26_7)*signed(FMAP_83_26);
			MULT_27(82)<=signed(DIN_27_7)*signed(FMAP_83_27);
			MULT_28(82)<=signed(DIN_28_7)*signed(FMAP_83_28);
			MULT_29(82)<=signed(DIN_29_7)*signed(FMAP_83_29);
			MULT_30(82)<=signed(DIN_30_7)*signed(FMAP_83_30);
			MULT_31(82)<=signed(DIN_31_7)*signed(FMAP_83_31);
			MULT_32(82)<=signed(DIN_32_7)*signed(FMAP_83_32);
			MULT_33(82)<=signed(DIN_33_7)*signed(FMAP_83_33);
			MULT_34(82)<=signed(DIN_34_7)*signed(FMAP_83_34);
			MULT_35(82)<=signed(DIN_35_7)*signed(FMAP_83_35);
			MULT_36(82)<=signed(DIN_36_7)*signed(FMAP_83_36);
			MULT_37(82)<=signed(DIN_37_7)*signed(FMAP_83_37);
			MULT_38(82)<=signed(DIN_38_7)*signed(FMAP_83_38);
			MULT_39(82)<=signed(DIN_39_7)*signed(FMAP_83_39);
			MULT_40(82)<=signed(DIN_40_7)*signed(FMAP_83_40);
			MULT_41(82)<=signed(DIN_41_7)*signed(FMAP_83_41);
			MULT_42(82)<=signed(DIN_42_7)*signed(FMAP_83_42);
			MULT_43(82)<=signed(DIN_43_7)*signed(FMAP_83_43);
			MULT_44(82)<=signed(DIN_44_7)*signed(FMAP_83_44);
			MULT_45(82)<=signed(DIN_45_7)*signed(FMAP_83_45);
			MULT_46(82)<=signed(DIN_46_7)*signed(FMAP_83_46);
			MULT_47(82)<=signed(DIN_47_7)*signed(FMAP_83_47);
			MULT_48(82)<=signed(DIN_48_7)*signed(FMAP_83_48);
			MULT_49(82)<=signed(DIN_49_7)*signed(FMAP_83_49);
			MULT_50(82)<=signed(DIN_50_7)*signed(FMAP_83_50);
			MULT_51(82)<=signed(DIN_51_7)*signed(FMAP_83_51);
			MULT_52(82)<=signed(DIN_52_7)*signed(FMAP_83_52);
			MULT_53(82)<=signed(DIN_53_7)*signed(FMAP_83_53);
			MULT_54(82)<=signed(DIN_54_7)*signed(FMAP_83_54);
			MULT_55(82)<=signed(DIN_55_7)*signed(FMAP_83_55);
			MULT_56(82)<=signed(DIN_56_7)*signed(FMAP_83_56);
			MULT_57(82)<=signed(DIN_57_7)*signed(FMAP_83_57);
			MULT_58(82)<=signed(DIN_58_7)*signed(FMAP_83_58);
			MULT_59(82)<=signed(DIN_59_7)*signed(FMAP_83_59);
			MULT_60(82)<=signed(DIN_60_7)*signed(FMAP_83_60);
			MULT_61(82)<=signed(DIN_61_7)*signed(FMAP_83_61);
			MULT_62(82)<=signed(DIN_62_7)*signed(FMAP_83_62);
			MULT_63(82)<=signed(DIN_63_7)*signed(FMAP_83_63);
			MULT_64(82)<=signed(DIN_64_7)*signed(FMAP_83_64);
			MULT_65(82)<=signed(DIN_65_7)*signed(FMAP_83_65);
			MULT_66(82)<=signed(DIN_66_7)*signed(FMAP_83_66);
			MULT_67(82)<=signed(DIN_67_7)*signed(FMAP_83_67);
			MULT_68(82)<=signed(DIN_68_7)*signed(FMAP_83_68);
			MULT_69(82)<=signed(DIN_69_7)*signed(FMAP_83_69);
			MULT_70(82)<=signed(DIN_70_7)*signed(FMAP_83_70);
			MULT_71(82)<=signed(DIN_71_7)*signed(FMAP_83_71);
			MULT_72(82)<=signed(DIN_72_7)*signed(FMAP_83_72);
			MULT_73(82)<=signed(DIN_73_7)*signed(FMAP_83_73);
			MULT_74(82)<=signed(DIN_74_7)*signed(FMAP_83_74);
			MULT_75(82)<=signed(DIN_75_7)*signed(FMAP_83_75);
			MULT_76(82)<=signed(DIN_76_7)*signed(FMAP_83_76);
			MULT_77(82)<=signed(DIN_77_7)*signed(FMAP_83_77);
			MULT_78(82)<=signed(DIN_78_7)*signed(FMAP_83_78);
			MULT_79(82)<=signed(DIN_79_7)*signed(FMAP_83_79);
			MULT_80(82)<=signed(DIN_80_7)*signed(FMAP_83_80);
			MULT_81(82)<=signed(DIN_81_7)*signed(FMAP_83_81);
			MULT_82(82)<=signed(DIN_82_7)*signed(FMAP_83_82);
			MULT_83(82)<=signed(DIN_83_7)*signed(FMAP_83_83);
			MULT_84(82)<=signed(DIN_84_7)*signed(FMAP_83_84);
			MULT_85(82)<=signed(DIN_85_7)*signed(FMAP_83_85);
			MULT_86(82)<=signed(DIN_86_7)*signed(FMAP_83_86);
			MULT_87(82)<=signed(DIN_87_7)*signed(FMAP_83_87);
			MULT_88(82)<=signed(DIN_88_7)*signed(FMAP_83_88);
			MULT_89(82)<=signed(DIN_89_7)*signed(FMAP_83_89);
			MULT_90(82)<=signed(DIN_90_7)*signed(FMAP_83_90);
			MULT_91(82)<=signed(DIN_91_7)*signed(FMAP_83_91);
			MULT_92(82)<=signed(DIN_92_7)*signed(FMAP_83_92);
			MULT_93(82)<=signed(DIN_93_7)*signed(FMAP_83_93);
			MULT_94(82)<=signed(DIN_94_7)*signed(FMAP_83_94);
			MULT_95(82)<=signed(DIN_95_7)*signed(FMAP_83_95);
			MULT_96(82)<=signed(DIN_96_7)*signed(FMAP_83_96);
			MULT_97(82)<=signed(DIN_97_7)*signed(FMAP_83_97);
			MULT_98(82)<=signed(DIN_98_7)*signed(FMAP_83_98);
			MULT_99(82)<=signed(DIN_99_7)*signed(FMAP_83_99);
			MULT_100(82)<=signed(DIN_100_7)*signed(FMAP_83_100);
			MULT_101(82)<=signed(DIN_101_7)*signed(FMAP_83_101);
			MULT_102(82)<=signed(DIN_102_7)*signed(FMAP_83_102);
			MULT_103(82)<=signed(DIN_103_7)*signed(FMAP_83_103);
			MULT_104(82)<=signed(DIN_104_7)*signed(FMAP_83_104);
			MULT_105(82)<=signed(DIN_105_7)*signed(FMAP_83_105);
			MULT_106(82)<=signed(DIN_106_7)*signed(FMAP_83_106);
			MULT_107(82)<=signed(DIN_107_7)*signed(FMAP_83_107);
			MULT_108(82)<=signed(DIN_108_7)*signed(FMAP_83_108);
			MULT_109(82)<=signed(DIN_109_7)*signed(FMAP_83_109);
			MULT_110(82)<=signed(DIN_110_7)*signed(FMAP_83_110);
			MULT_111(82)<=signed(DIN_111_7)*signed(FMAP_83_111);
			MULT_112(82)<=signed(DIN_112_7)*signed(FMAP_83_112);
			MULT_113(82)<=signed(DIN_113_7)*signed(FMAP_83_113);
			MULT_114(82)<=signed(DIN_114_7)*signed(FMAP_83_114);
			MULT_115(82)<=signed(DIN_115_7)*signed(FMAP_83_115);
			MULT_116(82)<=signed(DIN_116_7)*signed(FMAP_83_116);
			MULT_117(82)<=signed(DIN_117_7)*signed(FMAP_83_117);
			MULT_118(82)<=signed(DIN_118_7)*signed(FMAP_83_118);
			MULT_119(82)<=signed(DIN_119_7)*signed(FMAP_83_119);
			MULT_120(82)<=signed(DIN_120_7)*signed(FMAP_83_120);

			MULT_1(83)<=signed(DIN_1_7)*signed(FMAP_84_1);
			MULT_2(83)<=signed(DIN_2_7)*signed(FMAP_84_2);
			MULT_3(83)<=signed(DIN_3_7)*signed(FMAP_84_3);
			MULT_4(83)<=signed(DIN_4_7)*signed(FMAP_84_4);
			MULT_5(83)<=signed(DIN_5_7)*signed(FMAP_84_5);
			MULT_6(83)<=signed(DIN_6_7)*signed(FMAP_84_6);
			MULT_7(83)<=signed(DIN_7_7)*signed(FMAP_84_7);
			MULT_8(83)<=signed(DIN_8_7)*signed(FMAP_84_8);
			MULT_9(83)<=signed(DIN_9_7)*signed(FMAP_84_9);
			MULT_10(83)<=signed(DIN_10_7)*signed(FMAP_84_10);
			MULT_11(83)<=signed(DIN_11_7)*signed(FMAP_84_11);
			MULT_12(83)<=signed(DIN_12_7)*signed(FMAP_84_12);
			MULT_13(83)<=signed(DIN_13_7)*signed(FMAP_84_13);
			MULT_14(83)<=signed(DIN_14_7)*signed(FMAP_84_14);
			MULT_15(83)<=signed(DIN_15_7)*signed(FMAP_84_15);
			MULT_16(83)<=signed(DIN_16_7)*signed(FMAP_84_16);
			MULT_17(83)<=signed(DIN_17_7)*signed(FMAP_84_17);
			MULT_18(83)<=signed(DIN_18_7)*signed(FMAP_84_18);
			MULT_19(83)<=signed(DIN_19_7)*signed(FMAP_84_19);
			MULT_20(83)<=signed(DIN_20_7)*signed(FMAP_84_20);
			MULT_21(83)<=signed(DIN_21_7)*signed(FMAP_84_21);
			MULT_22(83)<=signed(DIN_22_7)*signed(FMAP_84_22);
			MULT_23(83)<=signed(DIN_23_7)*signed(FMAP_84_23);
			MULT_24(83)<=signed(DIN_24_7)*signed(FMAP_84_24);
			MULT_25(83)<=signed(DIN_25_7)*signed(FMAP_84_25);
			MULT_26(83)<=signed(DIN_26_7)*signed(FMAP_84_26);
			MULT_27(83)<=signed(DIN_27_7)*signed(FMAP_84_27);
			MULT_28(83)<=signed(DIN_28_7)*signed(FMAP_84_28);
			MULT_29(83)<=signed(DIN_29_7)*signed(FMAP_84_29);
			MULT_30(83)<=signed(DIN_30_7)*signed(FMAP_84_30);
			MULT_31(83)<=signed(DIN_31_7)*signed(FMAP_84_31);
			MULT_32(83)<=signed(DIN_32_7)*signed(FMAP_84_32);
			MULT_33(83)<=signed(DIN_33_7)*signed(FMAP_84_33);
			MULT_34(83)<=signed(DIN_34_7)*signed(FMAP_84_34);
			MULT_35(83)<=signed(DIN_35_7)*signed(FMAP_84_35);
			MULT_36(83)<=signed(DIN_36_7)*signed(FMAP_84_36);
			MULT_37(83)<=signed(DIN_37_7)*signed(FMAP_84_37);
			MULT_38(83)<=signed(DIN_38_7)*signed(FMAP_84_38);
			MULT_39(83)<=signed(DIN_39_7)*signed(FMAP_84_39);
			MULT_40(83)<=signed(DIN_40_7)*signed(FMAP_84_40);
			MULT_41(83)<=signed(DIN_41_7)*signed(FMAP_84_41);
			MULT_42(83)<=signed(DIN_42_7)*signed(FMAP_84_42);
			MULT_43(83)<=signed(DIN_43_7)*signed(FMAP_84_43);
			MULT_44(83)<=signed(DIN_44_7)*signed(FMAP_84_44);
			MULT_45(83)<=signed(DIN_45_7)*signed(FMAP_84_45);
			MULT_46(83)<=signed(DIN_46_7)*signed(FMAP_84_46);
			MULT_47(83)<=signed(DIN_47_7)*signed(FMAP_84_47);
			MULT_48(83)<=signed(DIN_48_7)*signed(FMAP_84_48);
			MULT_49(83)<=signed(DIN_49_7)*signed(FMAP_84_49);
			MULT_50(83)<=signed(DIN_50_7)*signed(FMAP_84_50);
			MULT_51(83)<=signed(DIN_51_7)*signed(FMAP_84_51);
			MULT_52(83)<=signed(DIN_52_7)*signed(FMAP_84_52);
			MULT_53(83)<=signed(DIN_53_7)*signed(FMAP_84_53);
			MULT_54(83)<=signed(DIN_54_7)*signed(FMAP_84_54);
			MULT_55(83)<=signed(DIN_55_7)*signed(FMAP_84_55);
			MULT_56(83)<=signed(DIN_56_7)*signed(FMAP_84_56);
			MULT_57(83)<=signed(DIN_57_7)*signed(FMAP_84_57);
			MULT_58(83)<=signed(DIN_58_7)*signed(FMAP_84_58);
			MULT_59(83)<=signed(DIN_59_7)*signed(FMAP_84_59);
			MULT_60(83)<=signed(DIN_60_7)*signed(FMAP_84_60);
			MULT_61(83)<=signed(DIN_61_7)*signed(FMAP_84_61);
			MULT_62(83)<=signed(DIN_62_7)*signed(FMAP_84_62);
			MULT_63(83)<=signed(DIN_63_7)*signed(FMAP_84_63);
			MULT_64(83)<=signed(DIN_64_7)*signed(FMAP_84_64);
			MULT_65(83)<=signed(DIN_65_7)*signed(FMAP_84_65);
			MULT_66(83)<=signed(DIN_66_7)*signed(FMAP_84_66);
			MULT_67(83)<=signed(DIN_67_7)*signed(FMAP_84_67);
			MULT_68(83)<=signed(DIN_68_7)*signed(FMAP_84_68);
			MULT_69(83)<=signed(DIN_69_7)*signed(FMAP_84_69);
			MULT_70(83)<=signed(DIN_70_7)*signed(FMAP_84_70);
			MULT_71(83)<=signed(DIN_71_7)*signed(FMAP_84_71);
			MULT_72(83)<=signed(DIN_72_7)*signed(FMAP_84_72);
			MULT_73(83)<=signed(DIN_73_7)*signed(FMAP_84_73);
			MULT_74(83)<=signed(DIN_74_7)*signed(FMAP_84_74);
			MULT_75(83)<=signed(DIN_75_7)*signed(FMAP_84_75);
			MULT_76(83)<=signed(DIN_76_7)*signed(FMAP_84_76);
			MULT_77(83)<=signed(DIN_77_7)*signed(FMAP_84_77);
			MULT_78(83)<=signed(DIN_78_7)*signed(FMAP_84_78);
			MULT_79(83)<=signed(DIN_79_7)*signed(FMAP_84_79);
			MULT_80(83)<=signed(DIN_80_7)*signed(FMAP_84_80);
			MULT_81(83)<=signed(DIN_81_7)*signed(FMAP_84_81);
			MULT_82(83)<=signed(DIN_82_7)*signed(FMAP_84_82);
			MULT_83(83)<=signed(DIN_83_7)*signed(FMAP_84_83);
			MULT_84(83)<=signed(DIN_84_7)*signed(FMAP_84_84);
			MULT_85(83)<=signed(DIN_85_7)*signed(FMAP_84_85);
			MULT_86(83)<=signed(DIN_86_7)*signed(FMAP_84_86);
			MULT_87(83)<=signed(DIN_87_7)*signed(FMAP_84_87);
			MULT_88(83)<=signed(DIN_88_7)*signed(FMAP_84_88);
			MULT_89(83)<=signed(DIN_89_7)*signed(FMAP_84_89);
			MULT_90(83)<=signed(DIN_90_7)*signed(FMAP_84_90);
			MULT_91(83)<=signed(DIN_91_7)*signed(FMAP_84_91);
			MULT_92(83)<=signed(DIN_92_7)*signed(FMAP_84_92);
			MULT_93(83)<=signed(DIN_93_7)*signed(FMAP_84_93);
			MULT_94(83)<=signed(DIN_94_7)*signed(FMAP_84_94);
			MULT_95(83)<=signed(DIN_95_7)*signed(FMAP_84_95);
			MULT_96(83)<=signed(DIN_96_7)*signed(FMAP_84_96);
			MULT_97(83)<=signed(DIN_97_7)*signed(FMAP_84_97);
			MULT_98(83)<=signed(DIN_98_7)*signed(FMAP_84_98);
			MULT_99(83)<=signed(DIN_99_7)*signed(FMAP_84_99);
			MULT_100(83)<=signed(DIN_100_7)*signed(FMAP_84_100);
			MULT_101(83)<=signed(DIN_101_7)*signed(FMAP_84_101);
			MULT_102(83)<=signed(DIN_102_7)*signed(FMAP_84_102);
			MULT_103(83)<=signed(DIN_103_7)*signed(FMAP_84_103);
			MULT_104(83)<=signed(DIN_104_7)*signed(FMAP_84_104);
			MULT_105(83)<=signed(DIN_105_7)*signed(FMAP_84_105);
			MULT_106(83)<=signed(DIN_106_7)*signed(FMAP_84_106);
			MULT_107(83)<=signed(DIN_107_7)*signed(FMAP_84_107);
			MULT_108(83)<=signed(DIN_108_7)*signed(FMAP_84_108);
			MULT_109(83)<=signed(DIN_109_7)*signed(FMAP_84_109);
			MULT_110(83)<=signed(DIN_110_7)*signed(FMAP_84_110);
			MULT_111(83)<=signed(DIN_111_7)*signed(FMAP_84_111);
			MULT_112(83)<=signed(DIN_112_7)*signed(FMAP_84_112);
			MULT_113(83)<=signed(DIN_113_7)*signed(FMAP_84_113);
			MULT_114(83)<=signed(DIN_114_7)*signed(FMAP_84_114);
			MULT_115(83)<=signed(DIN_115_7)*signed(FMAP_84_115);
			MULT_116(83)<=signed(DIN_116_7)*signed(FMAP_84_116);
			MULT_117(83)<=signed(DIN_117_7)*signed(FMAP_84_117);
			MULT_118(83)<=signed(DIN_118_7)*signed(FMAP_84_118);
			MULT_119(83)<=signed(DIN_119_7)*signed(FMAP_84_119);
			MULT_120(83)<=signed(DIN_120_7)*signed(FMAP_84_120);


                        EN_SUM_MULT_1<='1';

      -------------------------------------------- Enable MULT START --------------------------------------------				


		if EN_SUM_MULT_1 = '1' then
			------------------------------------STAGE-1--------------------------------------
			MULTS_1_1(0)<=signed(MULT_1(0)(MULT_SIZE-1) & MULT_1(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(0)(MULT_SIZE-1) & MULT_2(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(1)<=signed(MULT_1(1)(MULT_SIZE-1) & MULT_1(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(1)(MULT_SIZE-1) & MULT_2(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(2)<=signed(MULT_1(2)(MULT_SIZE-1) & MULT_1(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(2)(MULT_SIZE-1) & MULT_2(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(3)<=signed(MULT_1(3)(MULT_SIZE-1) & MULT_1(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(3)(MULT_SIZE-1) & MULT_2(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(4)<=signed(MULT_1(4)(MULT_SIZE-1) & MULT_1(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(4)(MULT_SIZE-1) & MULT_2(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(5)<=signed(MULT_1(5)(MULT_SIZE-1) & MULT_1(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(5)(MULT_SIZE-1) & MULT_2(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(6)<=signed(MULT_1(6)(MULT_SIZE-1) & MULT_1(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(6)(MULT_SIZE-1) & MULT_2(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(7)<=signed(MULT_1(7)(MULT_SIZE-1) & MULT_1(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(7)(MULT_SIZE-1) & MULT_2(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(8)<=signed(MULT_1(8)(MULT_SIZE-1) & MULT_1(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(8)(MULT_SIZE-1) & MULT_2(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(9)<=signed(MULT_1(9)(MULT_SIZE-1) & MULT_1(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(9)(MULT_SIZE-1) & MULT_2(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(10)<=signed(MULT_1(10)(MULT_SIZE-1) & MULT_1(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(10)(MULT_SIZE-1) & MULT_2(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(11)<=signed(MULT_1(11)(MULT_SIZE-1) & MULT_1(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(11)(MULT_SIZE-1) & MULT_2(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(12)<=signed(MULT_1(12)(MULT_SIZE-1) & MULT_1(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(12)(MULT_SIZE-1) & MULT_2(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(13)<=signed(MULT_1(13)(MULT_SIZE-1) & MULT_1(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(13)(MULT_SIZE-1) & MULT_2(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(14)<=signed(MULT_1(14)(MULT_SIZE-1) & MULT_1(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(14)(MULT_SIZE-1) & MULT_2(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(15)<=signed(MULT_1(15)(MULT_SIZE-1) & MULT_1(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(15)(MULT_SIZE-1) & MULT_2(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(16)<=signed(MULT_1(16)(MULT_SIZE-1) & MULT_1(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(16)(MULT_SIZE-1) & MULT_2(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(17)<=signed(MULT_1(17)(MULT_SIZE-1) & MULT_1(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(17)(MULT_SIZE-1) & MULT_2(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(18)<=signed(MULT_1(18)(MULT_SIZE-1) & MULT_1(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(18)(MULT_SIZE-1) & MULT_2(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(19)<=signed(MULT_1(19)(MULT_SIZE-1) & MULT_1(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(19)(MULT_SIZE-1) & MULT_2(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(20)<=signed(MULT_1(20)(MULT_SIZE-1) & MULT_1(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(20)(MULT_SIZE-1) & MULT_2(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(21)<=signed(MULT_1(21)(MULT_SIZE-1) & MULT_1(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(21)(MULT_SIZE-1) & MULT_2(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(22)<=signed(MULT_1(22)(MULT_SIZE-1) & MULT_1(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(22)(MULT_SIZE-1) & MULT_2(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(23)<=signed(MULT_1(23)(MULT_SIZE-1) & MULT_1(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(23)(MULT_SIZE-1) & MULT_2(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(24)<=signed(MULT_1(24)(MULT_SIZE-1) & MULT_1(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(24)(MULT_SIZE-1) & MULT_2(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(25)<=signed(MULT_1(25)(MULT_SIZE-1) & MULT_1(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(25)(MULT_SIZE-1) & MULT_2(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(26)<=signed(MULT_1(26)(MULT_SIZE-1) & MULT_1(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(26)(MULT_SIZE-1) & MULT_2(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(27)<=signed(MULT_1(27)(MULT_SIZE-1) & MULT_1(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(27)(MULT_SIZE-1) & MULT_2(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(28)<=signed(MULT_1(28)(MULT_SIZE-1) & MULT_1(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(28)(MULT_SIZE-1) & MULT_2(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(29)<=signed(MULT_1(29)(MULT_SIZE-1) & MULT_1(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(29)(MULT_SIZE-1) & MULT_2(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(30)<=signed(MULT_1(30)(MULT_SIZE-1) & MULT_1(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(30)(MULT_SIZE-1) & MULT_2(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(31)<=signed(MULT_1(31)(MULT_SIZE-1) & MULT_1(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(31)(MULT_SIZE-1) & MULT_2(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(32)<=signed(MULT_1(32)(MULT_SIZE-1) & MULT_1(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(32)(MULT_SIZE-1) & MULT_2(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(33)<=signed(MULT_1(33)(MULT_SIZE-1) & MULT_1(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(33)(MULT_SIZE-1) & MULT_2(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(34)<=signed(MULT_1(34)(MULT_SIZE-1) & MULT_1(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(34)(MULT_SIZE-1) & MULT_2(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(35)<=signed(MULT_1(35)(MULT_SIZE-1) & MULT_1(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(35)(MULT_SIZE-1) & MULT_2(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(36)<=signed(MULT_1(36)(MULT_SIZE-1) & MULT_1(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(36)(MULT_SIZE-1) & MULT_2(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(37)<=signed(MULT_1(37)(MULT_SIZE-1) & MULT_1(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(37)(MULT_SIZE-1) & MULT_2(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(38)<=signed(MULT_1(38)(MULT_SIZE-1) & MULT_1(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(38)(MULT_SIZE-1) & MULT_2(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(39)<=signed(MULT_1(39)(MULT_SIZE-1) & MULT_1(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(39)(MULT_SIZE-1) & MULT_2(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(40)<=signed(MULT_1(40)(MULT_SIZE-1) & MULT_1(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(40)(MULT_SIZE-1) & MULT_2(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(41)<=signed(MULT_1(41)(MULT_SIZE-1) & MULT_1(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(41)(MULT_SIZE-1) & MULT_2(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(42)<=signed(MULT_1(42)(MULT_SIZE-1) & MULT_1(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(42)(MULT_SIZE-1) & MULT_2(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(43)<=signed(MULT_1(43)(MULT_SIZE-1) & MULT_1(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(43)(MULT_SIZE-1) & MULT_2(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(44)<=signed(MULT_1(44)(MULT_SIZE-1) & MULT_1(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(44)(MULT_SIZE-1) & MULT_2(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(45)<=signed(MULT_1(45)(MULT_SIZE-1) & MULT_1(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(45)(MULT_SIZE-1) & MULT_2(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(46)<=signed(MULT_1(46)(MULT_SIZE-1) & MULT_1(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(46)(MULT_SIZE-1) & MULT_2(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(47)<=signed(MULT_1(47)(MULT_SIZE-1) & MULT_1(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(47)(MULT_SIZE-1) & MULT_2(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(48)<=signed(MULT_1(48)(MULT_SIZE-1) & MULT_1(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(48)(MULT_SIZE-1) & MULT_2(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(49)<=signed(MULT_1(49)(MULT_SIZE-1) & MULT_1(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(49)(MULT_SIZE-1) & MULT_2(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(50)<=signed(MULT_1(50)(MULT_SIZE-1) & MULT_1(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(50)(MULT_SIZE-1) & MULT_2(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(51)<=signed(MULT_1(51)(MULT_SIZE-1) & MULT_1(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(51)(MULT_SIZE-1) & MULT_2(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(52)<=signed(MULT_1(52)(MULT_SIZE-1) & MULT_1(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(52)(MULT_SIZE-1) & MULT_2(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(53)<=signed(MULT_1(53)(MULT_SIZE-1) & MULT_1(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(53)(MULT_SIZE-1) & MULT_2(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(54)<=signed(MULT_1(54)(MULT_SIZE-1) & MULT_1(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(54)(MULT_SIZE-1) & MULT_2(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(55)<=signed(MULT_1(55)(MULT_SIZE-1) & MULT_1(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(55)(MULT_SIZE-1) & MULT_2(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(56)<=signed(MULT_1(56)(MULT_SIZE-1) & MULT_1(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(56)(MULT_SIZE-1) & MULT_2(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(57)<=signed(MULT_1(57)(MULT_SIZE-1) & MULT_1(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(57)(MULT_SIZE-1) & MULT_2(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(58)<=signed(MULT_1(58)(MULT_SIZE-1) & MULT_1(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(58)(MULT_SIZE-1) & MULT_2(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(59)<=signed(MULT_1(59)(MULT_SIZE-1) & MULT_1(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(59)(MULT_SIZE-1) & MULT_2(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(60)<=signed(MULT_1(60)(MULT_SIZE-1) & MULT_1(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(60)(MULT_SIZE-1) & MULT_2(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(61)<=signed(MULT_1(61)(MULT_SIZE-1) & MULT_1(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(61)(MULT_SIZE-1) & MULT_2(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(62)<=signed(MULT_1(62)(MULT_SIZE-1) & MULT_1(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(62)(MULT_SIZE-1) & MULT_2(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(63)<=signed(MULT_1(63)(MULT_SIZE-1) & MULT_1(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(63)(MULT_SIZE-1) & MULT_2(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(64)<=signed(MULT_1(64)(MULT_SIZE-1) & MULT_1(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(64)(MULT_SIZE-1) & MULT_2(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(65)<=signed(MULT_1(65)(MULT_SIZE-1) & MULT_1(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(65)(MULT_SIZE-1) & MULT_2(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(66)<=signed(MULT_1(66)(MULT_SIZE-1) & MULT_1(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(66)(MULT_SIZE-1) & MULT_2(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(67)<=signed(MULT_1(67)(MULT_SIZE-1) & MULT_1(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(67)(MULT_SIZE-1) & MULT_2(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(68)<=signed(MULT_1(68)(MULT_SIZE-1) & MULT_1(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(68)(MULT_SIZE-1) & MULT_2(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(69)<=signed(MULT_1(69)(MULT_SIZE-1) & MULT_1(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(69)(MULT_SIZE-1) & MULT_2(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(70)<=signed(MULT_1(70)(MULT_SIZE-1) & MULT_1(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(70)(MULT_SIZE-1) & MULT_2(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(71)<=signed(MULT_1(71)(MULT_SIZE-1) & MULT_1(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(71)(MULT_SIZE-1) & MULT_2(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(72)<=signed(MULT_1(72)(MULT_SIZE-1) & MULT_1(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(72)(MULT_SIZE-1) & MULT_2(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(73)<=signed(MULT_1(73)(MULT_SIZE-1) & MULT_1(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(73)(MULT_SIZE-1) & MULT_2(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(74)<=signed(MULT_1(74)(MULT_SIZE-1) & MULT_1(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(74)(MULT_SIZE-1) & MULT_2(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(75)<=signed(MULT_1(75)(MULT_SIZE-1) & MULT_1(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(75)(MULT_SIZE-1) & MULT_2(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(76)<=signed(MULT_1(76)(MULT_SIZE-1) & MULT_1(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(76)(MULT_SIZE-1) & MULT_2(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(77)<=signed(MULT_1(77)(MULT_SIZE-1) & MULT_1(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(77)(MULT_SIZE-1) & MULT_2(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(78)<=signed(MULT_1(78)(MULT_SIZE-1) & MULT_1(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(78)(MULT_SIZE-1) & MULT_2(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(79)<=signed(MULT_1(79)(MULT_SIZE-1) & MULT_1(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(79)(MULT_SIZE-1) & MULT_2(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(80)<=signed(MULT_1(80)(MULT_SIZE-1) & MULT_1(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(80)(MULT_SIZE-1) & MULT_2(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(81)<=signed(MULT_1(81)(MULT_SIZE-1) & MULT_1(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(81)(MULT_SIZE-1) & MULT_2(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(82)<=signed(MULT_1(82)(MULT_SIZE-1) & MULT_1(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(82)(MULT_SIZE-1) & MULT_2(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1(83)<=signed(MULT_1(83)(MULT_SIZE-1) & MULT_1(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_2(83)(MULT_SIZE-1) & MULT_2(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_2(0)<=signed(MULT_3(0)(MULT_SIZE-1) & MULT_3(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(0)(MULT_SIZE-1) & MULT_4(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(1)<=signed(MULT_3(1)(MULT_SIZE-1) & MULT_3(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(1)(MULT_SIZE-1) & MULT_4(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(2)<=signed(MULT_3(2)(MULT_SIZE-1) & MULT_3(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(2)(MULT_SIZE-1) & MULT_4(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(3)<=signed(MULT_3(3)(MULT_SIZE-1) & MULT_3(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(3)(MULT_SIZE-1) & MULT_4(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(4)<=signed(MULT_3(4)(MULT_SIZE-1) & MULT_3(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(4)(MULT_SIZE-1) & MULT_4(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(5)<=signed(MULT_3(5)(MULT_SIZE-1) & MULT_3(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(5)(MULT_SIZE-1) & MULT_4(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(6)<=signed(MULT_3(6)(MULT_SIZE-1) & MULT_3(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(6)(MULT_SIZE-1) & MULT_4(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(7)<=signed(MULT_3(7)(MULT_SIZE-1) & MULT_3(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(7)(MULT_SIZE-1) & MULT_4(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(8)<=signed(MULT_3(8)(MULT_SIZE-1) & MULT_3(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(8)(MULT_SIZE-1) & MULT_4(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(9)<=signed(MULT_3(9)(MULT_SIZE-1) & MULT_3(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(9)(MULT_SIZE-1) & MULT_4(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(10)<=signed(MULT_3(10)(MULT_SIZE-1) & MULT_3(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(10)(MULT_SIZE-1) & MULT_4(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(11)<=signed(MULT_3(11)(MULT_SIZE-1) & MULT_3(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(11)(MULT_SIZE-1) & MULT_4(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(12)<=signed(MULT_3(12)(MULT_SIZE-1) & MULT_3(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(12)(MULT_SIZE-1) & MULT_4(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(13)<=signed(MULT_3(13)(MULT_SIZE-1) & MULT_3(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(13)(MULT_SIZE-1) & MULT_4(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(14)<=signed(MULT_3(14)(MULT_SIZE-1) & MULT_3(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(14)(MULT_SIZE-1) & MULT_4(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(15)<=signed(MULT_3(15)(MULT_SIZE-1) & MULT_3(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(15)(MULT_SIZE-1) & MULT_4(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(16)<=signed(MULT_3(16)(MULT_SIZE-1) & MULT_3(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(16)(MULT_SIZE-1) & MULT_4(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(17)<=signed(MULT_3(17)(MULT_SIZE-1) & MULT_3(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(17)(MULT_SIZE-1) & MULT_4(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(18)<=signed(MULT_3(18)(MULT_SIZE-1) & MULT_3(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(18)(MULT_SIZE-1) & MULT_4(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(19)<=signed(MULT_3(19)(MULT_SIZE-1) & MULT_3(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(19)(MULT_SIZE-1) & MULT_4(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(20)<=signed(MULT_3(20)(MULT_SIZE-1) & MULT_3(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(20)(MULT_SIZE-1) & MULT_4(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(21)<=signed(MULT_3(21)(MULT_SIZE-1) & MULT_3(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(21)(MULT_SIZE-1) & MULT_4(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(22)<=signed(MULT_3(22)(MULT_SIZE-1) & MULT_3(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(22)(MULT_SIZE-1) & MULT_4(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(23)<=signed(MULT_3(23)(MULT_SIZE-1) & MULT_3(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(23)(MULT_SIZE-1) & MULT_4(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(24)<=signed(MULT_3(24)(MULT_SIZE-1) & MULT_3(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(24)(MULT_SIZE-1) & MULT_4(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(25)<=signed(MULT_3(25)(MULT_SIZE-1) & MULT_3(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(25)(MULT_SIZE-1) & MULT_4(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(26)<=signed(MULT_3(26)(MULT_SIZE-1) & MULT_3(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(26)(MULT_SIZE-1) & MULT_4(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(27)<=signed(MULT_3(27)(MULT_SIZE-1) & MULT_3(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(27)(MULT_SIZE-1) & MULT_4(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(28)<=signed(MULT_3(28)(MULT_SIZE-1) & MULT_3(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(28)(MULT_SIZE-1) & MULT_4(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(29)<=signed(MULT_3(29)(MULT_SIZE-1) & MULT_3(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(29)(MULT_SIZE-1) & MULT_4(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(30)<=signed(MULT_3(30)(MULT_SIZE-1) & MULT_3(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(30)(MULT_SIZE-1) & MULT_4(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(31)<=signed(MULT_3(31)(MULT_SIZE-1) & MULT_3(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(31)(MULT_SIZE-1) & MULT_4(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(32)<=signed(MULT_3(32)(MULT_SIZE-1) & MULT_3(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(32)(MULT_SIZE-1) & MULT_4(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(33)<=signed(MULT_3(33)(MULT_SIZE-1) & MULT_3(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(33)(MULT_SIZE-1) & MULT_4(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(34)<=signed(MULT_3(34)(MULT_SIZE-1) & MULT_3(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(34)(MULT_SIZE-1) & MULT_4(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(35)<=signed(MULT_3(35)(MULT_SIZE-1) & MULT_3(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(35)(MULT_SIZE-1) & MULT_4(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(36)<=signed(MULT_3(36)(MULT_SIZE-1) & MULT_3(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(36)(MULT_SIZE-1) & MULT_4(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(37)<=signed(MULT_3(37)(MULT_SIZE-1) & MULT_3(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(37)(MULT_SIZE-1) & MULT_4(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(38)<=signed(MULT_3(38)(MULT_SIZE-1) & MULT_3(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(38)(MULT_SIZE-1) & MULT_4(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(39)<=signed(MULT_3(39)(MULT_SIZE-1) & MULT_3(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(39)(MULT_SIZE-1) & MULT_4(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(40)<=signed(MULT_3(40)(MULT_SIZE-1) & MULT_3(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(40)(MULT_SIZE-1) & MULT_4(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(41)<=signed(MULT_3(41)(MULT_SIZE-1) & MULT_3(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(41)(MULT_SIZE-1) & MULT_4(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(42)<=signed(MULT_3(42)(MULT_SIZE-1) & MULT_3(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(42)(MULT_SIZE-1) & MULT_4(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(43)<=signed(MULT_3(43)(MULT_SIZE-1) & MULT_3(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(43)(MULT_SIZE-1) & MULT_4(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(44)<=signed(MULT_3(44)(MULT_SIZE-1) & MULT_3(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(44)(MULT_SIZE-1) & MULT_4(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(45)<=signed(MULT_3(45)(MULT_SIZE-1) & MULT_3(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(45)(MULT_SIZE-1) & MULT_4(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(46)<=signed(MULT_3(46)(MULT_SIZE-1) & MULT_3(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(46)(MULT_SIZE-1) & MULT_4(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(47)<=signed(MULT_3(47)(MULT_SIZE-1) & MULT_3(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(47)(MULT_SIZE-1) & MULT_4(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(48)<=signed(MULT_3(48)(MULT_SIZE-1) & MULT_3(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(48)(MULT_SIZE-1) & MULT_4(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(49)<=signed(MULT_3(49)(MULT_SIZE-1) & MULT_3(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(49)(MULT_SIZE-1) & MULT_4(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(50)<=signed(MULT_3(50)(MULT_SIZE-1) & MULT_3(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(50)(MULT_SIZE-1) & MULT_4(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(51)<=signed(MULT_3(51)(MULT_SIZE-1) & MULT_3(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(51)(MULT_SIZE-1) & MULT_4(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(52)<=signed(MULT_3(52)(MULT_SIZE-1) & MULT_3(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(52)(MULT_SIZE-1) & MULT_4(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(53)<=signed(MULT_3(53)(MULT_SIZE-1) & MULT_3(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(53)(MULT_SIZE-1) & MULT_4(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(54)<=signed(MULT_3(54)(MULT_SIZE-1) & MULT_3(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(54)(MULT_SIZE-1) & MULT_4(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(55)<=signed(MULT_3(55)(MULT_SIZE-1) & MULT_3(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(55)(MULT_SIZE-1) & MULT_4(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(56)<=signed(MULT_3(56)(MULT_SIZE-1) & MULT_3(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(56)(MULT_SIZE-1) & MULT_4(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(57)<=signed(MULT_3(57)(MULT_SIZE-1) & MULT_3(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(57)(MULT_SIZE-1) & MULT_4(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(58)<=signed(MULT_3(58)(MULT_SIZE-1) & MULT_3(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(58)(MULT_SIZE-1) & MULT_4(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(59)<=signed(MULT_3(59)(MULT_SIZE-1) & MULT_3(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(59)(MULT_SIZE-1) & MULT_4(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(60)<=signed(MULT_3(60)(MULT_SIZE-1) & MULT_3(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(60)(MULT_SIZE-1) & MULT_4(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(61)<=signed(MULT_3(61)(MULT_SIZE-1) & MULT_3(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(61)(MULT_SIZE-1) & MULT_4(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(62)<=signed(MULT_3(62)(MULT_SIZE-1) & MULT_3(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(62)(MULT_SIZE-1) & MULT_4(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(63)<=signed(MULT_3(63)(MULT_SIZE-1) & MULT_3(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(63)(MULT_SIZE-1) & MULT_4(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(64)<=signed(MULT_3(64)(MULT_SIZE-1) & MULT_3(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(64)(MULT_SIZE-1) & MULT_4(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(65)<=signed(MULT_3(65)(MULT_SIZE-1) & MULT_3(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(65)(MULT_SIZE-1) & MULT_4(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(66)<=signed(MULT_3(66)(MULT_SIZE-1) & MULT_3(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(66)(MULT_SIZE-1) & MULT_4(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(67)<=signed(MULT_3(67)(MULT_SIZE-1) & MULT_3(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(67)(MULT_SIZE-1) & MULT_4(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(68)<=signed(MULT_3(68)(MULT_SIZE-1) & MULT_3(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(68)(MULT_SIZE-1) & MULT_4(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(69)<=signed(MULT_3(69)(MULT_SIZE-1) & MULT_3(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(69)(MULT_SIZE-1) & MULT_4(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(70)<=signed(MULT_3(70)(MULT_SIZE-1) & MULT_3(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(70)(MULT_SIZE-1) & MULT_4(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(71)<=signed(MULT_3(71)(MULT_SIZE-1) & MULT_3(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(71)(MULT_SIZE-1) & MULT_4(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(72)<=signed(MULT_3(72)(MULT_SIZE-1) & MULT_3(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(72)(MULT_SIZE-1) & MULT_4(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(73)<=signed(MULT_3(73)(MULT_SIZE-1) & MULT_3(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(73)(MULT_SIZE-1) & MULT_4(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(74)<=signed(MULT_3(74)(MULT_SIZE-1) & MULT_3(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(74)(MULT_SIZE-1) & MULT_4(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(75)<=signed(MULT_3(75)(MULT_SIZE-1) & MULT_3(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(75)(MULT_SIZE-1) & MULT_4(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(76)<=signed(MULT_3(76)(MULT_SIZE-1) & MULT_3(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(76)(MULT_SIZE-1) & MULT_4(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(77)<=signed(MULT_3(77)(MULT_SIZE-1) & MULT_3(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(77)(MULT_SIZE-1) & MULT_4(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(78)<=signed(MULT_3(78)(MULT_SIZE-1) & MULT_3(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(78)(MULT_SIZE-1) & MULT_4(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(79)<=signed(MULT_3(79)(MULT_SIZE-1) & MULT_3(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(79)(MULT_SIZE-1) & MULT_4(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(80)<=signed(MULT_3(80)(MULT_SIZE-1) & MULT_3(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(80)(MULT_SIZE-1) & MULT_4(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(81)<=signed(MULT_3(81)(MULT_SIZE-1) & MULT_3(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(81)(MULT_SIZE-1) & MULT_4(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(82)<=signed(MULT_3(82)(MULT_SIZE-1) & MULT_3(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(82)(MULT_SIZE-1) & MULT_4(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2(83)<=signed(MULT_3(83)(MULT_SIZE-1) & MULT_3(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_4(83)(MULT_SIZE-1) & MULT_4(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_3(0)<=signed(MULT_5(0)(MULT_SIZE-1) & MULT_5(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(0)(MULT_SIZE-1) & MULT_6(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(1)<=signed(MULT_5(1)(MULT_SIZE-1) & MULT_5(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(1)(MULT_SIZE-1) & MULT_6(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(2)<=signed(MULT_5(2)(MULT_SIZE-1) & MULT_5(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(2)(MULT_SIZE-1) & MULT_6(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(3)<=signed(MULT_5(3)(MULT_SIZE-1) & MULT_5(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(3)(MULT_SIZE-1) & MULT_6(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(4)<=signed(MULT_5(4)(MULT_SIZE-1) & MULT_5(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(4)(MULT_SIZE-1) & MULT_6(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(5)<=signed(MULT_5(5)(MULT_SIZE-1) & MULT_5(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(5)(MULT_SIZE-1) & MULT_6(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(6)<=signed(MULT_5(6)(MULT_SIZE-1) & MULT_5(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(6)(MULT_SIZE-1) & MULT_6(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(7)<=signed(MULT_5(7)(MULT_SIZE-1) & MULT_5(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(7)(MULT_SIZE-1) & MULT_6(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(8)<=signed(MULT_5(8)(MULT_SIZE-1) & MULT_5(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(8)(MULT_SIZE-1) & MULT_6(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(9)<=signed(MULT_5(9)(MULT_SIZE-1) & MULT_5(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(9)(MULT_SIZE-1) & MULT_6(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(10)<=signed(MULT_5(10)(MULT_SIZE-1) & MULT_5(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(10)(MULT_SIZE-1) & MULT_6(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(11)<=signed(MULT_5(11)(MULT_SIZE-1) & MULT_5(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(11)(MULT_SIZE-1) & MULT_6(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(12)<=signed(MULT_5(12)(MULT_SIZE-1) & MULT_5(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(12)(MULT_SIZE-1) & MULT_6(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(13)<=signed(MULT_5(13)(MULT_SIZE-1) & MULT_5(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(13)(MULT_SIZE-1) & MULT_6(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(14)<=signed(MULT_5(14)(MULT_SIZE-1) & MULT_5(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(14)(MULT_SIZE-1) & MULT_6(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(15)<=signed(MULT_5(15)(MULT_SIZE-1) & MULT_5(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(15)(MULT_SIZE-1) & MULT_6(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(16)<=signed(MULT_5(16)(MULT_SIZE-1) & MULT_5(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(16)(MULT_SIZE-1) & MULT_6(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(17)<=signed(MULT_5(17)(MULT_SIZE-1) & MULT_5(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(17)(MULT_SIZE-1) & MULT_6(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(18)<=signed(MULT_5(18)(MULT_SIZE-1) & MULT_5(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(18)(MULT_SIZE-1) & MULT_6(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(19)<=signed(MULT_5(19)(MULT_SIZE-1) & MULT_5(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(19)(MULT_SIZE-1) & MULT_6(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(20)<=signed(MULT_5(20)(MULT_SIZE-1) & MULT_5(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(20)(MULT_SIZE-1) & MULT_6(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(21)<=signed(MULT_5(21)(MULT_SIZE-1) & MULT_5(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(21)(MULT_SIZE-1) & MULT_6(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(22)<=signed(MULT_5(22)(MULT_SIZE-1) & MULT_5(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(22)(MULT_SIZE-1) & MULT_6(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(23)<=signed(MULT_5(23)(MULT_SIZE-1) & MULT_5(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(23)(MULT_SIZE-1) & MULT_6(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(24)<=signed(MULT_5(24)(MULT_SIZE-1) & MULT_5(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(24)(MULT_SIZE-1) & MULT_6(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(25)<=signed(MULT_5(25)(MULT_SIZE-1) & MULT_5(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(25)(MULT_SIZE-1) & MULT_6(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(26)<=signed(MULT_5(26)(MULT_SIZE-1) & MULT_5(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(26)(MULT_SIZE-1) & MULT_6(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(27)<=signed(MULT_5(27)(MULT_SIZE-1) & MULT_5(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(27)(MULT_SIZE-1) & MULT_6(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(28)<=signed(MULT_5(28)(MULT_SIZE-1) & MULT_5(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(28)(MULT_SIZE-1) & MULT_6(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(29)<=signed(MULT_5(29)(MULT_SIZE-1) & MULT_5(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(29)(MULT_SIZE-1) & MULT_6(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(30)<=signed(MULT_5(30)(MULT_SIZE-1) & MULT_5(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(30)(MULT_SIZE-1) & MULT_6(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(31)<=signed(MULT_5(31)(MULT_SIZE-1) & MULT_5(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(31)(MULT_SIZE-1) & MULT_6(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(32)<=signed(MULT_5(32)(MULT_SIZE-1) & MULT_5(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(32)(MULT_SIZE-1) & MULT_6(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(33)<=signed(MULT_5(33)(MULT_SIZE-1) & MULT_5(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(33)(MULT_SIZE-1) & MULT_6(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(34)<=signed(MULT_5(34)(MULT_SIZE-1) & MULT_5(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(34)(MULT_SIZE-1) & MULT_6(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(35)<=signed(MULT_5(35)(MULT_SIZE-1) & MULT_5(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(35)(MULT_SIZE-1) & MULT_6(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(36)<=signed(MULT_5(36)(MULT_SIZE-1) & MULT_5(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(36)(MULT_SIZE-1) & MULT_6(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(37)<=signed(MULT_5(37)(MULT_SIZE-1) & MULT_5(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(37)(MULT_SIZE-1) & MULT_6(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(38)<=signed(MULT_5(38)(MULT_SIZE-1) & MULT_5(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(38)(MULT_SIZE-1) & MULT_6(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(39)<=signed(MULT_5(39)(MULT_SIZE-1) & MULT_5(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(39)(MULT_SIZE-1) & MULT_6(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(40)<=signed(MULT_5(40)(MULT_SIZE-1) & MULT_5(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(40)(MULT_SIZE-1) & MULT_6(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(41)<=signed(MULT_5(41)(MULT_SIZE-1) & MULT_5(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(41)(MULT_SIZE-1) & MULT_6(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(42)<=signed(MULT_5(42)(MULT_SIZE-1) & MULT_5(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(42)(MULT_SIZE-1) & MULT_6(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(43)<=signed(MULT_5(43)(MULT_SIZE-1) & MULT_5(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(43)(MULT_SIZE-1) & MULT_6(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(44)<=signed(MULT_5(44)(MULT_SIZE-1) & MULT_5(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(44)(MULT_SIZE-1) & MULT_6(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(45)<=signed(MULT_5(45)(MULT_SIZE-1) & MULT_5(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(45)(MULT_SIZE-1) & MULT_6(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(46)<=signed(MULT_5(46)(MULT_SIZE-1) & MULT_5(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(46)(MULT_SIZE-1) & MULT_6(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(47)<=signed(MULT_5(47)(MULT_SIZE-1) & MULT_5(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(47)(MULT_SIZE-1) & MULT_6(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(48)<=signed(MULT_5(48)(MULT_SIZE-1) & MULT_5(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(48)(MULT_SIZE-1) & MULT_6(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(49)<=signed(MULT_5(49)(MULT_SIZE-1) & MULT_5(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(49)(MULT_SIZE-1) & MULT_6(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(50)<=signed(MULT_5(50)(MULT_SIZE-1) & MULT_5(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(50)(MULT_SIZE-1) & MULT_6(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(51)<=signed(MULT_5(51)(MULT_SIZE-1) & MULT_5(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(51)(MULT_SIZE-1) & MULT_6(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(52)<=signed(MULT_5(52)(MULT_SIZE-1) & MULT_5(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(52)(MULT_SIZE-1) & MULT_6(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(53)<=signed(MULT_5(53)(MULT_SIZE-1) & MULT_5(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(53)(MULT_SIZE-1) & MULT_6(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(54)<=signed(MULT_5(54)(MULT_SIZE-1) & MULT_5(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(54)(MULT_SIZE-1) & MULT_6(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(55)<=signed(MULT_5(55)(MULT_SIZE-1) & MULT_5(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(55)(MULT_SIZE-1) & MULT_6(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(56)<=signed(MULT_5(56)(MULT_SIZE-1) & MULT_5(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(56)(MULT_SIZE-1) & MULT_6(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(57)<=signed(MULT_5(57)(MULT_SIZE-1) & MULT_5(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(57)(MULT_SIZE-1) & MULT_6(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(58)<=signed(MULT_5(58)(MULT_SIZE-1) & MULT_5(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(58)(MULT_SIZE-1) & MULT_6(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(59)<=signed(MULT_5(59)(MULT_SIZE-1) & MULT_5(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(59)(MULT_SIZE-1) & MULT_6(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(60)<=signed(MULT_5(60)(MULT_SIZE-1) & MULT_5(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(60)(MULT_SIZE-1) & MULT_6(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(61)<=signed(MULT_5(61)(MULT_SIZE-1) & MULT_5(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(61)(MULT_SIZE-1) & MULT_6(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(62)<=signed(MULT_5(62)(MULT_SIZE-1) & MULT_5(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(62)(MULT_SIZE-1) & MULT_6(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(63)<=signed(MULT_5(63)(MULT_SIZE-1) & MULT_5(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(63)(MULT_SIZE-1) & MULT_6(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(64)<=signed(MULT_5(64)(MULT_SIZE-1) & MULT_5(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(64)(MULT_SIZE-1) & MULT_6(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(65)<=signed(MULT_5(65)(MULT_SIZE-1) & MULT_5(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(65)(MULT_SIZE-1) & MULT_6(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(66)<=signed(MULT_5(66)(MULT_SIZE-1) & MULT_5(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(66)(MULT_SIZE-1) & MULT_6(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(67)<=signed(MULT_5(67)(MULT_SIZE-1) & MULT_5(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(67)(MULT_SIZE-1) & MULT_6(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(68)<=signed(MULT_5(68)(MULT_SIZE-1) & MULT_5(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(68)(MULT_SIZE-1) & MULT_6(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(69)<=signed(MULT_5(69)(MULT_SIZE-1) & MULT_5(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(69)(MULT_SIZE-1) & MULT_6(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(70)<=signed(MULT_5(70)(MULT_SIZE-1) & MULT_5(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(70)(MULT_SIZE-1) & MULT_6(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(71)<=signed(MULT_5(71)(MULT_SIZE-1) & MULT_5(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(71)(MULT_SIZE-1) & MULT_6(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(72)<=signed(MULT_5(72)(MULT_SIZE-1) & MULT_5(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(72)(MULT_SIZE-1) & MULT_6(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(73)<=signed(MULT_5(73)(MULT_SIZE-1) & MULT_5(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(73)(MULT_SIZE-1) & MULT_6(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(74)<=signed(MULT_5(74)(MULT_SIZE-1) & MULT_5(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(74)(MULT_SIZE-1) & MULT_6(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(75)<=signed(MULT_5(75)(MULT_SIZE-1) & MULT_5(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(75)(MULT_SIZE-1) & MULT_6(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(76)<=signed(MULT_5(76)(MULT_SIZE-1) & MULT_5(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(76)(MULT_SIZE-1) & MULT_6(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(77)<=signed(MULT_5(77)(MULT_SIZE-1) & MULT_5(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(77)(MULT_SIZE-1) & MULT_6(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(78)<=signed(MULT_5(78)(MULT_SIZE-1) & MULT_5(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(78)(MULT_SIZE-1) & MULT_6(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(79)<=signed(MULT_5(79)(MULT_SIZE-1) & MULT_5(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(79)(MULT_SIZE-1) & MULT_6(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(80)<=signed(MULT_5(80)(MULT_SIZE-1) & MULT_5(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(80)(MULT_SIZE-1) & MULT_6(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(81)<=signed(MULT_5(81)(MULT_SIZE-1) & MULT_5(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(81)(MULT_SIZE-1) & MULT_6(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(82)<=signed(MULT_5(82)(MULT_SIZE-1) & MULT_5(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(82)(MULT_SIZE-1) & MULT_6(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3(83)<=signed(MULT_5(83)(MULT_SIZE-1) & MULT_5(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_6(83)(MULT_SIZE-1) & MULT_6(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_4(0)<=signed(MULT_7(0)(MULT_SIZE-1) & MULT_7(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(0)(MULT_SIZE-1) & MULT_8(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(1)<=signed(MULT_7(1)(MULT_SIZE-1) & MULT_7(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(1)(MULT_SIZE-1) & MULT_8(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(2)<=signed(MULT_7(2)(MULT_SIZE-1) & MULT_7(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(2)(MULT_SIZE-1) & MULT_8(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(3)<=signed(MULT_7(3)(MULT_SIZE-1) & MULT_7(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(3)(MULT_SIZE-1) & MULT_8(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(4)<=signed(MULT_7(4)(MULT_SIZE-1) & MULT_7(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(4)(MULT_SIZE-1) & MULT_8(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(5)<=signed(MULT_7(5)(MULT_SIZE-1) & MULT_7(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(5)(MULT_SIZE-1) & MULT_8(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(6)<=signed(MULT_7(6)(MULT_SIZE-1) & MULT_7(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(6)(MULT_SIZE-1) & MULT_8(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(7)<=signed(MULT_7(7)(MULT_SIZE-1) & MULT_7(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(7)(MULT_SIZE-1) & MULT_8(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(8)<=signed(MULT_7(8)(MULT_SIZE-1) & MULT_7(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(8)(MULT_SIZE-1) & MULT_8(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(9)<=signed(MULT_7(9)(MULT_SIZE-1) & MULT_7(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(9)(MULT_SIZE-1) & MULT_8(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(10)<=signed(MULT_7(10)(MULT_SIZE-1) & MULT_7(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(10)(MULT_SIZE-1) & MULT_8(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(11)<=signed(MULT_7(11)(MULT_SIZE-1) & MULT_7(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(11)(MULT_SIZE-1) & MULT_8(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(12)<=signed(MULT_7(12)(MULT_SIZE-1) & MULT_7(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(12)(MULT_SIZE-1) & MULT_8(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(13)<=signed(MULT_7(13)(MULT_SIZE-1) & MULT_7(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(13)(MULT_SIZE-1) & MULT_8(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(14)<=signed(MULT_7(14)(MULT_SIZE-1) & MULT_7(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(14)(MULT_SIZE-1) & MULT_8(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(15)<=signed(MULT_7(15)(MULT_SIZE-1) & MULT_7(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(15)(MULT_SIZE-1) & MULT_8(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(16)<=signed(MULT_7(16)(MULT_SIZE-1) & MULT_7(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(16)(MULT_SIZE-1) & MULT_8(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(17)<=signed(MULT_7(17)(MULT_SIZE-1) & MULT_7(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(17)(MULT_SIZE-1) & MULT_8(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(18)<=signed(MULT_7(18)(MULT_SIZE-1) & MULT_7(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(18)(MULT_SIZE-1) & MULT_8(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(19)<=signed(MULT_7(19)(MULT_SIZE-1) & MULT_7(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(19)(MULT_SIZE-1) & MULT_8(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(20)<=signed(MULT_7(20)(MULT_SIZE-1) & MULT_7(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(20)(MULT_SIZE-1) & MULT_8(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(21)<=signed(MULT_7(21)(MULT_SIZE-1) & MULT_7(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(21)(MULT_SIZE-1) & MULT_8(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(22)<=signed(MULT_7(22)(MULT_SIZE-1) & MULT_7(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(22)(MULT_SIZE-1) & MULT_8(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(23)<=signed(MULT_7(23)(MULT_SIZE-1) & MULT_7(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(23)(MULT_SIZE-1) & MULT_8(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(24)<=signed(MULT_7(24)(MULT_SIZE-1) & MULT_7(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(24)(MULT_SIZE-1) & MULT_8(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(25)<=signed(MULT_7(25)(MULT_SIZE-1) & MULT_7(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(25)(MULT_SIZE-1) & MULT_8(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(26)<=signed(MULT_7(26)(MULT_SIZE-1) & MULT_7(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(26)(MULT_SIZE-1) & MULT_8(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(27)<=signed(MULT_7(27)(MULT_SIZE-1) & MULT_7(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(27)(MULT_SIZE-1) & MULT_8(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(28)<=signed(MULT_7(28)(MULT_SIZE-1) & MULT_7(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(28)(MULT_SIZE-1) & MULT_8(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(29)<=signed(MULT_7(29)(MULT_SIZE-1) & MULT_7(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(29)(MULT_SIZE-1) & MULT_8(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(30)<=signed(MULT_7(30)(MULT_SIZE-1) & MULT_7(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(30)(MULT_SIZE-1) & MULT_8(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(31)<=signed(MULT_7(31)(MULT_SIZE-1) & MULT_7(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(31)(MULT_SIZE-1) & MULT_8(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(32)<=signed(MULT_7(32)(MULT_SIZE-1) & MULT_7(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(32)(MULT_SIZE-1) & MULT_8(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(33)<=signed(MULT_7(33)(MULT_SIZE-1) & MULT_7(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(33)(MULT_SIZE-1) & MULT_8(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(34)<=signed(MULT_7(34)(MULT_SIZE-1) & MULT_7(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(34)(MULT_SIZE-1) & MULT_8(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(35)<=signed(MULT_7(35)(MULT_SIZE-1) & MULT_7(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(35)(MULT_SIZE-1) & MULT_8(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(36)<=signed(MULT_7(36)(MULT_SIZE-1) & MULT_7(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(36)(MULT_SIZE-1) & MULT_8(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(37)<=signed(MULT_7(37)(MULT_SIZE-1) & MULT_7(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(37)(MULT_SIZE-1) & MULT_8(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(38)<=signed(MULT_7(38)(MULT_SIZE-1) & MULT_7(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(38)(MULT_SIZE-1) & MULT_8(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(39)<=signed(MULT_7(39)(MULT_SIZE-1) & MULT_7(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(39)(MULT_SIZE-1) & MULT_8(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(40)<=signed(MULT_7(40)(MULT_SIZE-1) & MULT_7(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(40)(MULT_SIZE-1) & MULT_8(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(41)<=signed(MULT_7(41)(MULT_SIZE-1) & MULT_7(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(41)(MULT_SIZE-1) & MULT_8(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(42)<=signed(MULT_7(42)(MULT_SIZE-1) & MULT_7(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(42)(MULT_SIZE-1) & MULT_8(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(43)<=signed(MULT_7(43)(MULT_SIZE-1) & MULT_7(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(43)(MULT_SIZE-1) & MULT_8(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(44)<=signed(MULT_7(44)(MULT_SIZE-1) & MULT_7(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(44)(MULT_SIZE-1) & MULT_8(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(45)<=signed(MULT_7(45)(MULT_SIZE-1) & MULT_7(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(45)(MULT_SIZE-1) & MULT_8(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(46)<=signed(MULT_7(46)(MULT_SIZE-1) & MULT_7(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(46)(MULT_SIZE-1) & MULT_8(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(47)<=signed(MULT_7(47)(MULT_SIZE-1) & MULT_7(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(47)(MULT_SIZE-1) & MULT_8(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(48)<=signed(MULT_7(48)(MULT_SIZE-1) & MULT_7(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(48)(MULT_SIZE-1) & MULT_8(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(49)<=signed(MULT_7(49)(MULT_SIZE-1) & MULT_7(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(49)(MULT_SIZE-1) & MULT_8(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(50)<=signed(MULT_7(50)(MULT_SIZE-1) & MULT_7(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(50)(MULT_SIZE-1) & MULT_8(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(51)<=signed(MULT_7(51)(MULT_SIZE-1) & MULT_7(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(51)(MULT_SIZE-1) & MULT_8(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(52)<=signed(MULT_7(52)(MULT_SIZE-1) & MULT_7(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(52)(MULT_SIZE-1) & MULT_8(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(53)<=signed(MULT_7(53)(MULT_SIZE-1) & MULT_7(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(53)(MULT_SIZE-1) & MULT_8(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(54)<=signed(MULT_7(54)(MULT_SIZE-1) & MULT_7(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(54)(MULT_SIZE-1) & MULT_8(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(55)<=signed(MULT_7(55)(MULT_SIZE-1) & MULT_7(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(55)(MULT_SIZE-1) & MULT_8(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(56)<=signed(MULT_7(56)(MULT_SIZE-1) & MULT_7(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(56)(MULT_SIZE-1) & MULT_8(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(57)<=signed(MULT_7(57)(MULT_SIZE-1) & MULT_7(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(57)(MULT_SIZE-1) & MULT_8(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(58)<=signed(MULT_7(58)(MULT_SIZE-1) & MULT_7(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(58)(MULT_SIZE-1) & MULT_8(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(59)<=signed(MULT_7(59)(MULT_SIZE-1) & MULT_7(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(59)(MULT_SIZE-1) & MULT_8(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(60)<=signed(MULT_7(60)(MULT_SIZE-1) & MULT_7(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(60)(MULT_SIZE-1) & MULT_8(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(61)<=signed(MULT_7(61)(MULT_SIZE-1) & MULT_7(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(61)(MULT_SIZE-1) & MULT_8(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(62)<=signed(MULT_7(62)(MULT_SIZE-1) & MULT_7(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(62)(MULT_SIZE-1) & MULT_8(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(63)<=signed(MULT_7(63)(MULT_SIZE-1) & MULT_7(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(63)(MULT_SIZE-1) & MULT_8(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(64)<=signed(MULT_7(64)(MULT_SIZE-1) & MULT_7(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(64)(MULT_SIZE-1) & MULT_8(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(65)<=signed(MULT_7(65)(MULT_SIZE-1) & MULT_7(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(65)(MULT_SIZE-1) & MULT_8(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(66)<=signed(MULT_7(66)(MULT_SIZE-1) & MULT_7(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(66)(MULT_SIZE-1) & MULT_8(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(67)<=signed(MULT_7(67)(MULT_SIZE-1) & MULT_7(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(67)(MULT_SIZE-1) & MULT_8(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(68)<=signed(MULT_7(68)(MULT_SIZE-1) & MULT_7(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(68)(MULT_SIZE-1) & MULT_8(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(69)<=signed(MULT_7(69)(MULT_SIZE-1) & MULT_7(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(69)(MULT_SIZE-1) & MULT_8(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(70)<=signed(MULT_7(70)(MULT_SIZE-1) & MULT_7(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(70)(MULT_SIZE-1) & MULT_8(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(71)<=signed(MULT_7(71)(MULT_SIZE-1) & MULT_7(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(71)(MULT_SIZE-1) & MULT_8(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(72)<=signed(MULT_7(72)(MULT_SIZE-1) & MULT_7(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(72)(MULT_SIZE-1) & MULT_8(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(73)<=signed(MULT_7(73)(MULT_SIZE-1) & MULT_7(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(73)(MULT_SIZE-1) & MULT_8(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(74)<=signed(MULT_7(74)(MULT_SIZE-1) & MULT_7(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(74)(MULT_SIZE-1) & MULT_8(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(75)<=signed(MULT_7(75)(MULT_SIZE-1) & MULT_7(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(75)(MULT_SIZE-1) & MULT_8(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(76)<=signed(MULT_7(76)(MULT_SIZE-1) & MULT_7(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(76)(MULT_SIZE-1) & MULT_8(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(77)<=signed(MULT_7(77)(MULT_SIZE-1) & MULT_7(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(77)(MULT_SIZE-1) & MULT_8(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(78)<=signed(MULT_7(78)(MULT_SIZE-1) & MULT_7(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(78)(MULT_SIZE-1) & MULT_8(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(79)<=signed(MULT_7(79)(MULT_SIZE-1) & MULT_7(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(79)(MULT_SIZE-1) & MULT_8(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(80)<=signed(MULT_7(80)(MULT_SIZE-1) & MULT_7(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(80)(MULT_SIZE-1) & MULT_8(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(81)<=signed(MULT_7(81)(MULT_SIZE-1) & MULT_7(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(81)(MULT_SIZE-1) & MULT_8(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(82)<=signed(MULT_7(82)(MULT_SIZE-1) & MULT_7(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(82)(MULT_SIZE-1) & MULT_8(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4(83)<=signed(MULT_7(83)(MULT_SIZE-1) & MULT_7(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_8(83)(MULT_SIZE-1) & MULT_8(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_5(0)<=signed(MULT_9(0)(MULT_SIZE-1) & MULT_9(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(0)(MULT_SIZE-1) & MULT_10(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(1)<=signed(MULT_9(1)(MULT_SIZE-1) & MULT_9(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(1)(MULT_SIZE-1) & MULT_10(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(2)<=signed(MULT_9(2)(MULT_SIZE-1) & MULT_9(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(2)(MULT_SIZE-1) & MULT_10(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(3)<=signed(MULT_9(3)(MULT_SIZE-1) & MULT_9(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(3)(MULT_SIZE-1) & MULT_10(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(4)<=signed(MULT_9(4)(MULT_SIZE-1) & MULT_9(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(4)(MULT_SIZE-1) & MULT_10(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(5)<=signed(MULT_9(5)(MULT_SIZE-1) & MULT_9(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(5)(MULT_SIZE-1) & MULT_10(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(6)<=signed(MULT_9(6)(MULT_SIZE-1) & MULT_9(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(6)(MULT_SIZE-1) & MULT_10(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(7)<=signed(MULT_9(7)(MULT_SIZE-1) & MULT_9(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(7)(MULT_SIZE-1) & MULT_10(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(8)<=signed(MULT_9(8)(MULT_SIZE-1) & MULT_9(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(8)(MULT_SIZE-1) & MULT_10(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(9)<=signed(MULT_9(9)(MULT_SIZE-1) & MULT_9(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(9)(MULT_SIZE-1) & MULT_10(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(10)<=signed(MULT_9(10)(MULT_SIZE-1) & MULT_9(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(10)(MULT_SIZE-1) & MULT_10(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(11)<=signed(MULT_9(11)(MULT_SIZE-1) & MULT_9(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(11)(MULT_SIZE-1) & MULT_10(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(12)<=signed(MULT_9(12)(MULT_SIZE-1) & MULT_9(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(12)(MULT_SIZE-1) & MULT_10(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(13)<=signed(MULT_9(13)(MULT_SIZE-1) & MULT_9(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(13)(MULT_SIZE-1) & MULT_10(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(14)<=signed(MULT_9(14)(MULT_SIZE-1) & MULT_9(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(14)(MULT_SIZE-1) & MULT_10(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(15)<=signed(MULT_9(15)(MULT_SIZE-1) & MULT_9(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(15)(MULT_SIZE-1) & MULT_10(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(16)<=signed(MULT_9(16)(MULT_SIZE-1) & MULT_9(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(16)(MULT_SIZE-1) & MULT_10(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(17)<=signed(MULT_9(17)(MULT_SIZE-1) & MULT_9(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(17)(MULT_SIZE-1) & MULT_10(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(18)<=signed(MULT_9(18)(MULT_SIZE-1) & MULT_9(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(18)(MULT_SIZE-1) & MULT_10(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(19)<=signed(MULT_9(19)(MULT_SIZE-1) & MULT_9(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(19)(MULT_SIZE-1) & MULT_10(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(20)<=signed(MULT_9(20)(MULT_SIZE-1) & MULT_9(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(20)(MULT_SIZE-1) & MULT_10(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(21)<=signed(MULT_9(21)(MULT_SIZE-1) & MULT_9(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(21)(MULT_SIZE-1) & MULT_10(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(22)<=signed(MULT_9(22)(MULT_SIZE-1) & MULT_9(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(22)(MULT_SIZE-1) & MULT_10(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(23)<=signed(MULT_9(23)(MULT_SIZE-1) & MULT_9(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(23)(MULT_SIZE-1) & MULT_10(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(24)<=signed(MULT_9(24)(MULT_SIZE-1) & MULT_9(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(24)(MULT_SIZE-1) & MULT_10(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(25)<=signed(MULT_9(25)(MULT_SIZE-1) & MULT_9(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(25)(MULT_SIZE-1) & MULT_10(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(26)<=signed(MULT_9(26)(MULT_SIZE-1) & MULT_9(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(26)(MULT_SIZE-1) & MULT_10(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(27)<=signed(MULT_9(27)(MULT_SIZE-1) & MULT_9(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(27)(MULT_SIZE-1) & MULT_10(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(28)<=signed(MULT_9(28)(MULT_SIZE-1) & MULT_9(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(28)(MULT_SIZE-1) & MULT_10(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(29)<=signed(MULT_9(29)(MULT_SIZE-1) & MULT_9(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(29)(MULT_SIZE-1) & MULT_10(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(30)<=signed(MULT_9(30)(MULT_SIZE-1) & MULT_9(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(30)(MULT_SIZE-1) & MULT_10(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(31)<=signed(MULT_9(31)(MULT_SIZE-1) & MULT_9(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(31)(MULT_SIZE-1) & MULT_10(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(32)<=signed(MULT_9(32)(MULT_SIZE-1) & MULT_9(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(32)(MULT_SIZE-1) & MULT_10(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(33)<=signed(MULT_9(33)(MULT_SIZE-1) & MULT_9(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(33)(MULT_SIZE-1) & MULT_10(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(34)<=signed(MULT_9(34)(MULT_SIZE-1) & MULT_9(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(34)(MULT_SIZE-1) & MULT_10(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(35)<=signed(MULT_9(35)(MULT_SIZE-1) & MULT_9(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(35)(MULT_SIZE-1) & MULT_10(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(36)<=signed(MULT_9(36)(MULT_SIZE-1) & MULT_9(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(36)(MULT_SIZE-1) & MULT_10(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(37)<=signed(MULT_9(37)(MULT_SIZE-1) & MULT_9(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(37)(MULT_SIZE-1) & MULT_10(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(38)<=signed(MULT_9(38)(MULT_SIZE-1) & MULT_9(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(38)(MULT_SIZE-1) & MULT_10(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(39)<=signed(MULT_9(39)(MULT_SIZE-1) & MULT_9(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(39)(MULT_SIZE-1) & MULT_10(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(40)<=signed(MULT_9(40)(MULT_SIZE-1) & MULT_9(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(40)(MULT_SIZE-1) & MULT_10(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(41)<=signed(MULT_9(41)(MULT_SIZE-1) & MULT_9(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(41)(MULT_SIZE-1) & MULT_10(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(42)<=signed(MULT_9(42)(MULT_SIZE-1) & MULT_9(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(42)(MULT_SIZE-1) & MULT_10(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(43)<=signed(MULT_9(43)(MULT_SIZE-1) & MULT_9(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(43)(MULT_SIZE-1) & MULT_10(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(44)<=signed(MULT_9(44)(MULT_SIZE-1) & MULT_9(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(44)(MULT_SIZE-1) & MULT_10(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(45)<=signed(MULT_9(45)(MULT_SIZE-1) & MULT_9(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(45)(MULT_SIZE-1) & MULT_10(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(46)<=signed(MULT_9(46)(MULT_SIZE-1) & MULT_9(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(46)(MULT_SIZE-1) & MULT_10(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(47)<=signed(MULT_9(47)(MULT_SIZE-1) & MULT_9(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(47)(MULT_SIZE-1) & MULT_10(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(48)<=signed(MULT_9(48)(MULT_SIZE-1) & MULT_9(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(48)(MULT_SIZE-1) & MULT_10(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(49)<=signed(MULT_9(49)(MULT_SIZE-1) & MULT_9(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(49)(MULT_SIZE-1) & MULT_10(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(50)<=signed(MULT_9(50)(MULT_SIZE-1) & MULT_9(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(50)(MULT_SIZE-1) & MULT_10(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(51)<=signed(MULT_9(51)(MULT_SIZE-1) & MULT_9(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(51)(MULT_SIZE-1) & MULT_10(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(52)<=signed(MULT_9(52)(MULT_SIZE-1) & MULT_9(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(52)(MULT_SIZE-1) & MULT_10(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(53)<=signed(MULT_9(53)(MULT_SIZE-1) & MULT_9(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(53)(MULT_SIZE-1) & MULT_10(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(54)<=signed(MULT_9(54)(MULT_SIZE-1) & MULT_9(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(54)(MULT_SIZE-1) & MULT_10(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(55)<=signed(MULT_9(55)(MULT_SIZE-1) & MULT_9(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(55)(MULT_SIZE-1) & MULT_10(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(56)<=signed(MULT_9(56)(MULT_SIZE-1) & MULT_9(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(56)(MULT_SIZE-1) & MULT_10(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(57)<=signed(MULT_9(57)(MULT_SIZE-1) & MULT_9(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(57)(MULT_SIZE-1) & MULT_10(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(58)<=signed(MULT_9(58)(MULT_SIZE-1) & MULT_9(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(58)(MULT_SIZE-1) & MULT_10(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(59)<=signed(MULT_9(59)(MULT_SIZE-1) & MULT_9(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(59)(MULT_SIZE-1) & MULT_10(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(60)<=signed(MULT_9(60)(MULT_SIZE-1) & MULT_9(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(60)(MULT_SIZE-1) & MULT_10(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(61)<=signed(MULT_9(61)(MULT_SIZE-1) & MULT_9(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(61)(MULT_SIZE-1) & MULT_10(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(62)<=signed(MULT_9(62)(MULT_SIZE-1) & MULT_9(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(62)(MULT_SIZE-1) & MULT_10(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(63)<=signed(MULT_9(63)(MULT_SIZE-1) & MULT_9(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(63)(MULT_SIZE-1) & MULT_10(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(64)<=signed(MULT_9(64)(MULT_SIZE-1) & MULT_9(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(64)(MULT_SIZE-1) & MULT_10(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(65)<=signed(MULT_9(65)(MULT_SIZE-1) & MULT_9(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(65)(MULT_SIZE-1) & MULT_10(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(66)<=signed(MULT_9(66)(MULT_SIZE-1) & MULT_9(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(66)(MULT_SIZE-1) & MULT_10(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(67)<=signed(MULT_9(67)(MULT_SIZE-1) & MULT_9(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(67)(MULT_SIZE-1) & MULT_10(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(68)<=signed(MULT_9(68)(MULT_SIZE-1) & MULT_9(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(68)(MULT_SIZE-1) & MULT_10(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(69)<=signed(MULT_9(69)(MULT_SIZE-1) & MULT_9(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(69)(MULT_SIZE-1) & MULT_10(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(70)<=signed(MULT_9(70)(MULT_SIZE-1) & MULT_9(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(70)(MULT_SIZE-1) & MULT_10(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(71)<=signed(MULT_9(71)(MULT_SIZE-1) & MULT_9(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(71)(MULT_SIZE-1) & MULT_10(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(72)<=signed(MULT_9(72)(MULT_SIZE-1) & MULT_9(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(72)(MULT_SIZE-1) & MULT_10(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(73)<=signed(MULT_9(73)(MULT_SIZE-1) & MULT_9(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(73)(MULT_SIZE-1) & MULT_10(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(74)<=signed(MULT_9(74)(MULT_SIZE-1) & MULT_9(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(74)(MULT_SIZE-1) & MULT_10(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(75)<=signed(MULT_9(75)(MULT_SIZE-1) & MULT_9(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(75)(MULT_SIZE-1) & MULT_10(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(76)<=signed(MULT_9(76)(MULT_SIZE-1) & MULT_9(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(76)(MULT_SIZE-1) & MULT_10(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(77)<=signed(MULT_9(77)(MULT_SIZE-1) & MULT_9(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(77)(MULT_SIZE-1) & MULT_10(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(78)<=signed(MULT_9(78)(MULT_SIZE-1) & MULT_9(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(78)(MULT_SIZE-1) & MULT_10(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(79)<=signed(MULT_9(79)(MULT_SIZE-1) & MULT_9(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(79)(MULT_SIZE-1) & MULT_10(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(80)<=signed(MULT_9(80)(MULT_SIZE-1) & MULT_9(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(80)(MULT_SIZE-1) & MULT_10(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(81)<=signed(MULT_9(81)(MULT_SIZE-1) & MULT_9(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(81)(MULT_SIZE-1) & MULT_10(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(82)<=signed(MULT_9(82)(MULT_SIZE-1) & MULT_9(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(82)(MULT_SIZE-1) & MULT_10(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5(83)<=signed(MULT_9(83)(MULT_SIZE-1) & MULT_9(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_10(83)(MULT_SIZE-1) & MULT_10(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_6(0)<=signed(MULT_11(0)(MULT_SIZE-1) & MULT_11(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(0)(MULT_SIZE-1) & MULT_12(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(1)<=signed(MULT_11(1)(MULT_SIZE-1) & MULT_11(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(1)(MULT_SIZE-1) & MULT_12(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(2)<=signed(MULT_11(2)(MULT_SIZE-1) & MULT_11(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(2)(MULT_SIZE-1) & MULT_12(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(3)<=signed(MULT_11(3)(MULT_SIZE-1) & MULT_11(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(3)(MULT_SIZE-1) & MULT_12(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(4)<=signed(MULT_11(4)(MULT_SIZE-1) & MULT_11(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(4)(MULT_SIZE-1) & MULT_12(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(5)<=signed(MULT_11(5)(MULT_SIZE-1) & MULT_11(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(5)(MULT_SIZE-1) & MULT_12(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(6)<=signed(MULT_11(6)(MULT_SIZE-1) & MULT_11(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(6)(MULT_SIZE-1) & MULT_12(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(7)<=signed(MULT_11(7)(MULT_SIZE-1) & MULT_11(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(7)(MULT_SIZE-1) & MULT_12(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(8)<=signed(MULT_11(8)(MULT_SIZE-1) & MULT_11(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(8)(MULT_SIZE-1) & MULT_12(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(9)<=signed(MULT_11(9)(MULT_SIZE-1) & MULT_11(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(9)(MULT_SIZE-1) & MULT_12(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(10)<=signed(MULT_11(10)(MULT_SIZE-1) & MULT_11(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(10)(MULT_SIZE-1) & MULT_12(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(11)<=signed(MULT_11(11)(MULT_SIZE-1) & MULT_11(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(11)(MULT_SIZE-1) & MULT_12(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(12)<=signed(MULT_11(12)(MULT_SIZE-1) & MULT_11(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(12)(MULT_SIZE-1) & MULT_12(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(13)<=signed(MULT_11(13)(MULT_SIZE-1) & MULT_11(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(13)(MULT_SIZE-1) & MULT_12(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(14)<=signed(MULT_11(14)(MULT_SIZE-1) & MULT_11(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(14)(MULT_SIZE-1) & MULT_12(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(15)<=signed(MULT_11(15)(MULT_SIZE-1) & MULT_11(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(15)(MULT_SIZE-1) & MULT_12(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(16)<=signed(MULT_11(16)(MULT_SIZE-1) & MULT_11(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(16)(MULT_SIZE-1) & MULT_12(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(17)<=signed(MULT_11(17)(MULT_SIZE-1) & MULT_11(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(17)(MULT_SIZE-1) & MULT_12(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(18)<=signed(MULT_11(18)(MULT_SIZE-1) & MULT_11(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(18)(MULT_SIZE-1) & MULT_12(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(19)<=signed(MULT_11(19)(MULT_SIZE-1) & MULT_11(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(19)(MULT_SIZE-1) & MULT_12(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(20)<=signed(MULT_11(20)(MULT_SIZE-1) & MULT_11(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(20)(MULT_SIZE-1) & MULT_12(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(21)<=signed(MULT_11(21)(MULT_SIZE-1) & MULT_11(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(21)(MULT_SIZE-1) & MULT_12(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(22)<=signed(MULT_11(22)(MULT_SIZE-1) & MULT_11(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(22)(MULT_SIZE-1) & MULT_12(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(23)<=signed(MULT_11(23)(MULT_SIZE-1) & MULT_11(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(23)(MULT_SIZE-1) & MULT_12(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(24)<=signed(MULT_11(24)(MULT_SIZE-1) & MULT_11(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(24)(MULT_SIZE-1) & MULT_12(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(25)<=signed(MULT_11(25)(MULT_SIZE-1) & MULT_11(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(25)(MULT_SIZE-1) & MULT_12(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(26)<=signed(MULT_11(26)(MULT_SIZE-1) & MULT_11(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(26)(MULT_SIZE-1) & MULT_12(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(27)<=signed(MULT_11(27)(MULT_SIZE-1) & MULT_11(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(27)(MULT_SIZE-1) & MULT_12(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(28)<=signed(MULT_11(28)(MULT_SIZE-1) & MULT_11(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(28)(MULT_SIZE-1) & MULT_12(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(29)<=signed(MULT_11(29)(MULT_SIZE-1) & MULT_11(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(29)(MULT_SIZE-1) & MULT_12(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(30)<=signed(MULT_11(30)(MULT_SIZE-1) & MULT_11(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(30)(MULT_SIZE-1) & MULT_12(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(31)<=signed(MULT_11(31)(MULT_SIZE-1) & MULT_11(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(31)(MULT_SIZE-1) & MULT_12(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(32)<=signed(MULT_11(32)(MULT_SIZE-1) & MULT_11(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(32)(MULT_SIZE-1) & MULT_12(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(33)<=signed(MULT_11(33)(MULT_SIZE-1) & MULT_11(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(33)(MULT_SIZE-1) & MULT_12(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(34)<=signed(MULT_11(34)(MULT_SIZE-1) & MULT_11(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(34)(MULT_SIZE-1) & MULT_12(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(35)<=signed(MULT_11(35)(MULT_SIZE-1) & MULT_11(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(35)(MULT_SIZE-1) & MULT_12(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(36)<=signed(MULT_11(36)(MULT_SIZE-1) & MULT_11(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(36)(MULT_SIZE-1) & MULT_12(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(37)<=signed(MULT_11(37)(MULT_SIZE-1) & MULT_11(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(37)(MULT_SIZE-1) & MULT_12(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(38)<=signed(MULT_11(38)(MULT_SIZE-1) & MULT_11(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(38)(MULT_SIZE-1) & MULT_12(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(39)<=signed(MULT_11(39)(MULT_SIZE-1) & MULT_11(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(39)(MULT_SIZE-1) & MULT_12(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(40)<=signed(MULT_11(40)(MULT_SIZE-1) & MULT_11(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(40)(MULT_SIZE-1) & MULT_12(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(41)<=signed(MULT_11(41)(MULT_SIZE-1) & MULT_11(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(41)(MULT_SIZE-1) & MULT_12(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(42)<=signed(MULT_11(42)(MULT_SIZE-1) & MULT_11(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(42)(MULT_SIZE-1) & MULT_12(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(43)<=signed(MULT_11(43)(MULT_SIZE-1) & MULT_11(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(43)(MULT_SIZE-1) & MULT_12(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(44)<=signed(MULT_11(44)(MULT_SIZE-1) & MULT_11(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(44)(MULT_SIZE-1) & MULT_12(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(45)<=signed(MULT_11(45)(MULT_SIZE-1) & MULT_11(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(45)(MULT_SIZE-1) & MULT_12(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(46)<=signed(MULT_11(46)(MULT_SIZE-1) & MULT_11(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(46)(MULT_SIZE-1) & MULT_12(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(47)<=signed(MULT_11(47)(MULT_SIZE-1) & MULT_11(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(47)(MULT_SIZE-1) & MULT_12(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(48)<=signed(MULT_11(48)(MULT_SIZE-1) & MULT_11(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(48)(MULT_SIZE-1) & MULT_12(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(49)<=signed(MULT_11(49)(MULT_SIZE-1) & MULT_11(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(49)(MULT_SIZE-1) & MULT_12(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(50)<=signed(MULT_11(50)(MULT_SIZE-1) & MULT_11(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(50)(MULT_SIZE-1) & MULT_12(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(51)<=signed(MULT_11(51)(MULT_SIZE-1) & MULT_11(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(51)(MULT_SIZE-1) & MULT_12(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(52)<=signed(MULT_11(52)(MULT_SIZE-1) & MULT_11(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(52)(MULT_SIZE-1) & MULT_12(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(53)<=signed(MULT_11(53)(MULT_SIZE-1) & MULT_11(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(53)(MULT_SIZE-1) & MULT_12(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(54)<=signed(MULT_11(54)(MULT_SIZE-1) & MULT_11(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(54)(MULT_SIZE-1) & MULT_12(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(55)<=signed(MULT_11(55)(MULT_SIZE-1) & MULT_11(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(55)(MULT_SIZE-1) & MULT_12(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(56)<=signed(MULT_11(56)(MULT_SIZE-1) & MULT_11(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(56)(MULT_SIZE-1) & MULT_12(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(57)<=signed(MULT_11(57)(MULT_SIZE-1) & MULT_11(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(57)(MULT_SIZE-1) & MULT_12(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(58)<=signed(MULT_11(58)(MULT_SIZE-1) & MULT_11(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(58)(MULT_SIZE-1) & MULT_12(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(59)<=signed(MULT_11(59)(MULT_SIZE-1) & MULT_11(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(59)(MULT_SIZE-1) & MULT_12(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(60)<=signed(MULT_11(60)(MULT_SIZE-1) & MULT_11(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(60)(MULT_SIZE-1) & MULT_12(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(61)<=signed(MULT_11(61)(MULT_SIZE-1) & MULT_11(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(61)(MULT_SIZE-1) & MULT_12(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(62)<=signed(MULT_11(62)(MULT_SIZE-1) & MULT_11(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(62)(MULT_SIZE-1) & MULT_12(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(63)<=signed(MULT_11(63)(MULT_SIZE-1) & MULT_11(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(63)(MULT_SIZE-1) & MULT_12(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(64)<=signed(MULT_11(64)(MULT_SIZE-1) & MULT_11(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(64)(MULT_SIZE-1) & MULT_12(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(65)<=signed(MULT_11(65)(MULT_SIZE-1) & MULT_11(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(65)(MULT_SIZE-1) & MULT_12(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(66)<=signed(MULT_11(66)(MULT_SIZE-1) & MULT_11(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(66)(MULT_SIZE-1) & MULT_12(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(67)<=signed(MULT_11(67)(MULT_SIZE-1) & MULT_11(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(67)(MULT_SIZE-1) & MULT_12(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(68)<=signed(MULT_11(68)(MULT_SIZE-1) & MULT_11(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(68)(MULT_SIZE-1) & MULT_12(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(69)<=signed(MULT_11(69)(MULT_SIZE-1) & MULT_11(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(69)(MULT_SIZE-1) & MULT_12(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(70)<=signed(MULT_11(70)(MULT_SIZE-1) & MULT_11(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(70)(MULT_SIZE-1) & MULT_12(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(71)<=signed(MULT_11(71)(MULT_SIZE-1) & MULT_11(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(71)(MULT_SIZE-1) & MULT_12(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(72)<=signed(MULT_11(72)(MULT_SIZE-1) & MULT_11(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(72)(MULT_SIZE-1) & MULT_12(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(73)<=signed(MULT_11(73)(MULT_SIZE-1) & MULT_11(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(73)(MULT_SIZE-1) & MULT_12(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(74)<=signed(MULT_11(74)(MULT_SIZE-1) & MULT_11(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(74)(MULT_SIZE-1) & MULT_12(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(75)<=signed(MULT_11(75)(MULT_SIZE-1) & MULT_11(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(75)(MULT_SIZE-1) & MULT_12(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(76)<=signed(MULT_11(76)(MULT_SIZE-1) & MULT_11(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(76)(MULT_SIZE-1) & MULT_12(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(77)<=signed(MULT_11(77)(MULT_SIZE-1) & MULT_11(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(77)(MULT_SIZE-1) & MULT_12(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(78)<=signed(MULT_11(78)(MULT_SIZE-1) & MULT_11(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(78)(MULT_SIZE-1) & MULT_12(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(79)<=signed(MULT_11(79)(MULT_SIZE-1) & MULT_11(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(79)(MULT_SIZE-1) & MULT_12(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(80)<=signed(MULT_11(80)(MULT_SIZE-1) & MULT_11(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(80)(MULT_SIZE-1) & MULT_12(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(81)<=signed(MULT_11(81)(MULT_SIZE-1) & MULT_11(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(81)(MULT_SIZE-1) & MULT_12(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(82)<=signed(MULT_11(82)(MULT_SIZE-1) & MULT_11(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(82)(MULT_SIZE-1) & MULT_12(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6(83)<=signed(MULT_11(83)(MULT_SIZE-1) & MULT_11(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_12(83)(MULT_SIZE-1) & MULT_12(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_7(0)<=signed(MULT_13(0)(MULT_SIZE-1) & MULT_13(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(0)(MULT_SIZE-1) & MULT_14(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(1)<=signed(MULT_13(1)(MULT_SIZE-1) & MULT_13(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(1)(MULT_SIZE-1) & MULT_14(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(2)<=signed(MULT_13(2)(MULT_SIZE-1) & MULT_13(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(2)(MULT_SIZE-1) & MULT_14(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(3)<=signed(MULT_13(3)(MULT_SIZE-1) & MULT_13(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(3)(MULT_SIZE-1) & MULT_14(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(4)<=signed(MULT_13(4)(MULT_SIZE-1) & MULT_13(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(4)(MULT_SIZE-1) & MULT_14(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(5)<=signed(MULT_13(5)(MULT_SIZE-1) & MULT_13(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(5)(MULT_SIZE-1) & MULT_14(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(6)<=signed(MULT_13(6)(MULT_SIZE-1) & MULT_13(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(6)(MULT_SIZE-1) & MULT_14(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(7)<=signed(MULT_13(7)(MULT_SIZE-1) & MULT_13(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(7)(MULT_SIZE-1) & MULT_14(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(8)<=signed(MULT_13(8)(MULT_SIZE-1) & MULT_13(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(8)(MULT_SIZE-1) & MULT_14(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(9)<=signed(MULT_13(9)(MULT_SIZE-1) & MULT_13(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(9)(MULT_SIZE-1) & MULT_14(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(10)<=signed(MULT_13(10)(MULT_SIZE-1) & MULT_13(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(10)(MULT_SIZE-1) & MULT_14(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(11)<=signed(MULT_13(11)(MULT_SIZE-1) & MULT_13(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(11)(MULT_SIZE-1) & MULT_14(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(12)<=signed(MULT_13(12)(MULT_SIZE-1) & MULT_13(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(12)(MULT_SIZE-1) & MULT_14(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(13)<=signed(MULT_13(13)(MULT_SIZE-1) & MULT_13(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(13)(MULT_SIZE-1) & MULT_14(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(14)<=signed(MULT_13(14)(MULT_SIZE-1) & MULT_13(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(14)(MULT_SIZE-1) & MULT_14(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(15)<=signed(MULT_13(15)(MULT_SIZE-1) & MULT_13(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(15)(MULT_SIZE-1) & MULT_14(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(16)<=signed(MULT_13(16)(MULT_SIZE-1) & MULT_13(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(16)(MULT_SIZE-1) & MULT_14(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(17)<=signed(MULT_13(17)(MULT_SIZE-1) & MULT_13(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(17)(MULT_SIZE-1) & MULT_14(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(18)<=signed(MULT_13(18)(MULT_SIZE-1) & MULT_13(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(18)(MULT_SIZE-1) & MULT_14(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(19)<=signed(MULT_13(19)(MULT_SIZE-1) & MULT_13(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(19)(MULT_SIZE-1) & MULT_14(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(20)<=signed(MULT_13(20)(MULT_SIZE-1) & MULT_13(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(20)(MULT_SIZE-1) & MULT_14(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(21)<=signed(MULT_13(21)(MULT_SIZE-1) & MULT_13(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(21)(MULT_SIZE-1) & MULT_14(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(22)<=signed(MULT_13(22)(MULT_SIZE-1) & MULT_13(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(22)(MULT_SIZE-1) & MULT_14(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(23)<=signed(MULT_13(23)(MULT_SIZE-1) & MULT_13(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(23)(MULT_SIZE-1) & MULT_14(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(24)<=signed(MULT_13(24)(MULT_SIZE-1) & MULT_13(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(24)(MULT_SIZE-1) & MULT_14(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(25)<=signed(MULT_13(25)(MULT_SIZE-1) & MULT_13(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(25)(MULT_SIZE-1) & MULT_14(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(26)<=signed(MULT_13(26)(MULT_SIZE-1) & MULT_13(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(26)(MULT_SIZE-1) & MULT_14(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(27)<=signed(MULT_13(27)(MULT_SIZE-1) & MULT_13(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(27)(MULT_SIZE-1) & MULT_14(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(28)<=signed(MULT_13(28)(MULT_SIZE-1) & MULT_13(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(28)(MULT_SIZE-1) & MULT_14(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(29)<=signed(MULT_13(29)(MULT_SIZE-1) & MULT_13(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(29)(MULT_SIZE-1) & MULT_14(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(30)<=signed(MULT_13(30)(MULT_SIZE-1) & MULT_13(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(30)(MULT_SIZE-1) & MULT_14(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(31)<=signed(MULT_13(31)(MULT_SIZE-1) & MULT_13(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(31)(MULT_SIZE-1) & MULT_14(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(32)<=signed(MULT_13(32)(MULT_SIZE-1) & MULT_13(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(32)(MULT_SIZE-1) & MULT_14(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(33)<=signed(MULT_13(33)(MULT_SIZE-1) & MULT_13(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(33)(MULT_SIZE-1) & MULT_14(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(34)<=signed(MULT_13(34)(MULT_SIZE-1) & MULT_13(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(34)(MULT_SIZE-1) & MULT_14(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(35)<=signed(MULT_13(35)(MULT_SIZE-1) & MULT_13(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(35)(MULT_SIZE-1) & MULT_14(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(36)<=signed(MULT_13(36)(MULT_SIZE-1) & MULT_13(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(36)(MULT_SIZE-1) & MULT_14(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(37)<=signed(MULT_13(37)(MULT_SIZE-1) & MULT_13(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(37)(MULT_SIZE-1) & MULT_14(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(38)<=signed(MULT_13(38)(MULT_SIZE-1) & MULT_13(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(38)(MULT_SIZE-1) & MULT_14(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(39)<=signed(MULT_13(39)(MULT_SIZE-1) & MULT_13(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(39)(MULT_SIZE-1) & MULT_14(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(40)<=signed(MULT_13(40)(MULT_SIZE-1) & MULT_13(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(40)(MULT_SIZE-1) & MULT_14(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(41)<=signed(MULT_13(41)(MULT_SIZE-1) & MULT_13(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(41)(MULT_SIZE-1) & MULT_14(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(42)<=signed(MULT_13(42)(MULT_SIZE-1) & MULT_13(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(42)(MULT_SIZE-1) & MULT_14(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(43)<=signed(MULT_13(43)(MULT_SIZE-1) & MULT_13(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(43)(MULT_SIZE-1) & MULT_14(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(44)<=signed(MULT_13(44)(MULT_SIZE-1) & MULT_13(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(44)(MULT_SIZE-1) & MULT_14(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(45)<=signed(MULT_13(45)(MULT_SIZE-1) & MULT_13(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(45)(MULT_SIZE-1) & MULT_14(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(46)<=signed(MULT_13(46)(MULT_SIZE-1) & MULT_13(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(46)(MULT_SIZE-1) & MULT_14(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(47)<=signed(MULT_13(47)(MULT_SIZE-1) & MULT_13(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(47)(MULT_SIZE-1) & MULT_14(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(48)<=signed(MULT_13(48)(MULT_SIZE-1) & MULT_13(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(48)(MULT_SIZE-1) & MULT_14(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(49)<=signed(MULT_13(49)(MULT_SIZE-1) & MULT_13(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(49)(MULT_SIZE-1) & MULT_14(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(50)<=signed(MULT_13(50)(MULT_SIZE-1) & MULT_13(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(50)(MULT_SIZE-1) & MULT_14(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(51)<=signed(MULT_13(51)(MULT_SIZE-1) & MULT_13(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(51)(MULT_SIZE-1) & MULT_14(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(52)<=signed(MULT_13(52)(MULT_SIZE-1) & MULT_13(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(52)(MULT_SIZE-1) & MULT_14(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(53)<=signed(MULT_13(53)(MULT_SIZE-1) & MULT_13(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(53)(MULT_SIZE-1) & MULT_14(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(54)<=signed(MULT_13(54)(MULT_SIZE-1) & MULT_13(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(54)(MULT_SIZE-1) & MULT_14(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(55)<=signed(MULT_13(55)(MULT_SIZE-1) & MULT_13(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(55)(MULT_SIZE-1) & MULT_14(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(56)<=signed(MULT_13(56)(MULT_SIZE-1) & MULT_13(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(56)(MULT_SIZE-1) & MULT_14(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(57)<=signed(MULT_13(57)(MULT_SIZE-1) & MULT_13(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(57)(MULT_SIZE-1) & MULT_14(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(58)<=signed(MULT_13(58)(MULT_SIZE-1) & MULT_13(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(58)(MULT_SIZE-1) & MULT_14(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(59)<=signed(MULT_13(59)(MULT_SIZE-1) & MULT_13(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(59)(MULT_SIZE-1) & MULT_14(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(60)<=signed(MULT_13(60)(MULT_SIZE-1) & MULT_13(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(60)(MULT_SIZE-1) & MULT_14(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(61)<=signed(MULT_13(61)(MULT_SIZE-1) & MULT_13(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(61)(MULT_SIZE-1) & MULT_14(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(62)<=signed(MULT_13(62)(MULT_SIZE-1) & MULT_13(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(62)(MULT_SIZE-1) & MULT_14(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(63)<=signed(MULT_13(63)(MULT_SIZE-1) & MULT_13(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(63)(MULT_SIZE-1) & MULT_14(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(64)<=signed(MULT_13(64)(MULT_SIZE-1) & MULT_13(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(64)(MULT_SIZE-1) & MULT_14(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(65)<=signed(MULT_13(65)(MULT_SIZE-1) & MULT_13(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(65)(MULT_SIZE-1) & MULT_14(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(66)<=signed(MULT_13(66)(MULT_SIZE-1) & MULT_13(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(66)(MULT_SIZE-1) & MULT_14(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(67)<=signed(MULT_13(67)(MULT_SIZE-1) & MULT_13(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(67)(MULT_SIZE-1) & MULT_14(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(68)<=signed(MULT_13(68)(MULT_SIZE-1) & MULT_13(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(68)(MULT_SIZE-1) & MULT_14(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(69)<=signed(MULT_13(69)(MULT_SIZE-1) & MULT_13(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(69)(MULT_SIZE-1) & MULT_14(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(70)<=signed(MULT_13(70)(MULT_SIZE-1) & MULT_13(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(70)(MULT_SIZE-1) & MULT_14(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(71)<=signed(MULT_13(71)(MULT_SIZE-1) & MULT_13(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(71)(MULT_SIZE-1) & MULT_14(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(72)<=signed(MULT_13(72)(MULT_SIZE-1) & MULT_13(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(72)(MULT_SIZE-1) & MULT_14(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(73)<=signed(MULT_13(73)(MULT_SIZE-1) & MULT_13(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(73)(MULT_SIZE-1) & MULT_14(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(74)<=signed(MULT_13(74)(MULT_SIZE-1) & MULT_13(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(74)(MULT_SIZE-1) & MULT_14(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(75)<=signed(MULT_13(75)(MULT_SIZE-1) & MULT_13(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(75)(MULT_SIZE-1) & MULT_14(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(76)<=signed(MULT_13(76)(MULT_SIZE-1) & MULT_13(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(76)(MULT_SIZE-1) & MULT_14(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(77)<=signed(MULT_13(77)(MULT_SIZE-1) & MULT_13(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(77)(MULT_SIZE-1) & MULT_14(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(78)<=signed(MULT_13(78)(MULT_SIZE-1) & MULT_13(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(78)(MULT_SIZE-1) & MULT_14(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(79)<=signed(MULT_13(79)(MULT_SIZE-1) & MULT_13(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(79)(MULT_SIZE-1) & MULT_14(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(80)<=signed(MULT_13(80)(MULT_SIZE-1) & MULT_13(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(80)(MULT_SIZE-1) & MULT_14(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(81)<=signed(MULT_13(81)(MULT_SIZE-1) & MULT_13(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(81)(MULT_SIZE-1) & MULT_14(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(82)<=signed(MULT_13(82)(MULT_SIZE-1) & MULT_13(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(82)(MULT_SIZE-1) & MULT_14(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7(83)<=signed(MULT_13(83)(MULT_SIZE-1) & MULT_13(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_14(83)(MULT_SIZE-1) & MULT_14(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_8(0)<=signed(MULT_15(0)(MULT_SIZE-1) & MULT_15(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(0)(MULT_SIZE-1) & MULT_16(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(1)<=signed(MULT_15(1)(MULT_SIZE-1) & MULT_15(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(1)(MULT_SIZE-1) & MULT_16(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(2)<=signed(MULT_15(2)(MULT_SIZE-1) & MULT_15(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(2)(MULT_SIZE-1) & MULT_16(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(3)<=signed(MULT_15(3)(MULT_SIZE-1) & MULT_15(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(3)(MULT_SIZE-1) & MULT_16(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(4)<=signed(MULT_15(4)(MULT_SIZE-1) & MULT_15(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(4)(MULT_SIZE-1) & MULT_16(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(5)<=signed(MULT_15(5)(MULT_SIZE-1) & MULT_15(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(5)(MULT_SIZE-1) & MULT_16(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(6)<=signed(MULT_15(6)(MULT_SIZE-1) & MULT_15(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(6)(MULT_SIZE-1) & MULT_16(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(7)<=signed(MULT_15(7)(MULT_SIZE-1) & MULT_15(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(7)(MULT_SIZE-1) & MULT_16(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(8)<=signed(MULT_15(8)(MULT_SIZE-1) & MULT_15(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(8)(MULT_SIZE-1) & MULT_16(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(9)<=signed(MULT_15(9)(MULT_SIZE-1) & MULT_15(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(9)(MULT_SIZE-1) & MULT_16(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(10)<=signed(MULT_15(10)(MULT_SIZE-1) & MULT_15(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(10)(MULT_SIZE-1) & MULT_16(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(11)<=signed(MULT_15(11)(MULT_SIZE-1) & MULT_15(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(11)(MULT_SIZE-1) & MULT_16(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(12)<=signed(MULT_15(12)(MULT_SIZE-1) & MULT_15(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(12)(MULT_SIZE-1) & MULT_16(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(13)<=signed(MULT_15(13)(MULT_SIZE-1) & MULT_15(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(13)(MULT_SIZE-1) & MULT_16(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(14)<=signed(MULT_15(14)(MULT_SIZE-1) & MULT_15(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(14)(MULT_SIZE-1) & MULT_16(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(15)<=signed(MULT_15(15)(MULT_SIZE-1) & MULT_15(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(15)(MULT_SIZE-1) & MULT_16(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(16)<=signed(MULT_15(16)(MULT_SIZE-1) & MULT_15(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(16)(MULT_SIZE-1) & MULT_16(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(17)<=signed(MULT_15(17)(MULT_SIZE-1) & MULT_15(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(17)(MULT_SIZE-1) & MULT_16(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(18)<=signed(MULT_15(18)(MULT_SIZE-1) & MULT_15(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(18)(MULT_SIZE-1) & MULT_16(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(19)<=signed(MULT_15(19)(MULT_SIZE-1) & MULT_15(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(19)(MULT_SIZE-1) & MULT_16(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(20)<=signed(MULT_15(20)(MULT_SIZE-1) & MULT_15(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(20)(MULT_SIZE-1) & MULT_16(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(21)<=signed(MULT_15(21)(MULT_SIZE-1) & MULT_15(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(21)(MULT_SIZE-1) & MULT_16(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(22)<=signed(MULT_15(22)(MULT_SIZE-1) & MULT_15(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(22)(MULT_SIZE-1) & MULT_16(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(23)<=signed(MULT_15(23)(MULT_SIZE-1) & MULT_15(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(23)(MULT_SIZE-1) & MULT_16(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(24)<=signed(MULT_15(24)(MULT_SIZE-1) & MULT_15(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(24)(MULT_SIZE-1) & MULT_16(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(25)<=signed(MULT_15(25)(MULT_SIZE-1) & MULT_15(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(25)(MULT_SIZE-1) & MULT_16(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(26)<=signed(MULT_15(26)(MULT_SIZE-1) & MULT_15(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(26)(MULT_SIZE-1) & MULT_16(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(27)<=signed(MULT_15(27)(MULT_SIZE-1) & MULT_15(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(27)(MULT_SIZE-1) & MULT_16(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(28)<=signed(MULT_15(28)(MULT_SIZE-1) & MULT_15(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(28)(MULT_SIZE-1) & MULT_16(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(29)<=signed(MULT_15(29)(MULT_SIZE-1) & MULT_15(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(29)(MULT_SIZE-1) & MULT_16(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(30)<=signed(MULT_15(30)(MULT_SIZE-1) & MULT_15(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(30)(MULT_SIZE-1) & MULT_16(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(31)<=signed(MULT_15(31)(MULT_SIZE-1) & MULT_15(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(31)(MULT_SIZE-1) & MULT_16(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(32)<=signed(MULT_15(32)(MULT_SIZE-1) & MULT_15(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(32)(MULT_SIZE-1) & MULT_16(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(33)<=signed(MULT_15(33)(MULT_SIZE-1) & MULT_15(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(33)(MULT_SIZE-1) & MULT_16(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(34)<=signed(MULT_15(34)(MULT_SIZE-1) & MULT_15(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(34)(MULT_SIZE-1) & MULT_16(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(35)<=signed(MULT_15(35)(MULT_SIZE-1) & MULT_15(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(35)(MULT_SIZE-1) & MULT_16(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(36)<=signed(MULT_15(36)(MULT_SIZE-1) & MULT_15(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(36)(MULT_SIZE-1) & MULT_16(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(37)<=signed(MULT_15(37)(MULT_SIZE-1) & MULT_15(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(37)(MULT_SIZE-1) & MULT_16(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(38)<=signed(MULT_15(38)(MULT_SIZE-1) & MULT_15(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(38)(MULT_SIZE-1) & MULT_16(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(39)<=signed(MULT_15(39)(MULT_SIZE-1) & MULT_15(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(39)(MULT_SIZE-1) & MULT_16(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(40)<=signed(MULT_15(40)(MULT_SIZE-1) & MULT_15(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(40)(MULT_SIZE-1) & MULT_16(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(41)<=signed(MULT_15(41)(MULT_SIZE-1) & MULT_15(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(41)(MULT_SIZE-1) & MULT_16(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(42)<=signed(MULT_15(42)(MULT_SIZE-1) & MULT_15(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(42)(MULT_SIZE-1) & MULT_16(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(43)<=signed(MULT_15(43)(MULT_SIZE-1) & MULT_15(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(43)(MULT_SIZE-1) & MULT_16(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(44)<=signed(MULT_15(44)(MULT_SIZE-1) & MULT_15(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(44)(MULT_SIZE-1) & MULT_16(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(45)<=signed(MULT_15(45)(MULT_SIZE-1) & MULT_15(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(45)(MULT_SIZE-1) & MULT_16(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(46)<=signed(MULT_15(46)(MULT_SIZE-1) & MULT_15(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(46)(MULT_SIZE-1) & MULT_16(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(47)<=signed(MULT_15(47)(MULT_SIZE-1) & MULT_15(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(47)(MULT_SIZE-1) & MULT_16(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(48)<=signed(MULT_15(48)(MULT_SIZE-1) & MULT_15(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(48)(MULT_SIZE-1) & MULT_16(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(49)<=signed(MULT_15(49)(MULT_SIZE-1) & MULT_15(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(49)(MULT_SIZE-1) & MULT_16(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(50)<=signed(MULT_15(50)(MULT_SIZE-1) & MULT_15(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(50)(MULT_SIZE-1) & MULT_16(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(51)<=signed(MULT_15(51)(MULT_SIZE-1) & MULT_15(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(51)(MULT_SIZE-1) & MULT_16(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(52)<=signed(MULT_15(52)(MULT_SIZE-1) & MULT_15(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(52)(MULT_SIZE-1) & MULT_16(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(53)<=signed(MULT_15(53)(MULT_SIZE-1) & MULT_15(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(53)(MULT_SIZE-1) & MULT_16(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(54)<=signed(MULT_15(54)(MULT_SIZE-1) & MULT_15(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(54)(MULT_SIZE-1) & MULT_16(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(55)<=signed(MULT_15(55)(MULT_SIZE-1) & MULT_15(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(55)(MULT_SIZE-1) & MULT_16(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(56)<=signed(MULT_15(56)(MULT_SIZE-1) & MULT_15(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(56)(MULT_SIZE-1) & MULT_16(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(57)<=signed(MULT_15(57)(MULT_SIZE-1) & MULT_15(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(57)(MULT_SIZE-1) & MULT_16(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(58)<=signed(MULT_15(58)(MULT_SIZE-1) & MULT_15(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(58)(MULT_SIZE-1) & MULT_16(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(59)<=signed(MULT_15(59)(MULT_SIZE-1) & MULT_15(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(59)(MULT_SIZE-1) & MULT_16(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(60)<=signed(MULT_15(60)(MULT_SIZE-1) & MULT_15(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(60)(MULT_SIZE-1) & MULT_16(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(61)<=signed(MULT_15(61)(MULT_SIZE-1) & MULT_15(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(61)(MULT_SIZE-1) & MULT_16(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(62)<=signed(MULT_15(62)(MULT_SIZE-1) & MULT_15(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(62)(MULT_SIZE-1) & MULT_16(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(63)<=signed(MULT_15(63)(MULT_SIZE-1) & MULT_15(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(63)(MULT_SIZE-1) & MULT_16(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(64)<=signed(MULT_15(64)(MULT_SIZE-1) & MULT_15(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(64)(MULT_SIZE-1) & MULT_16(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(65)<=signed(MULT_15(65)(MULT_SIZE-1) & MULT_15(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(65)(MULT_SIZE-1) & MULT_16(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(66)<=signed(MULT_15(66)(MULT_SIZE-1) & MULT_15(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(66)(MULT_SIZE-1) & MULT_16(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(67)<=signed(MULT_15(67)(MULT_SIZE-1) & MULT_15(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(67)(MULT_SIZE-1) & MULT_16(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(68)<=signed(MULT_15(68)(MULT_SIZE-1) & MULT_15(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(68)(MULT_SIZE-1) & MULT_16(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(69)<=signed(MULT_15(69)(MULT_SIZE-1) & MULT_15(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(69)(MULT_SIZE-1) & MULT_16(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(70)<=signed(MULT_15(70)(MULT_SIZE-1) & MULT_15(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(70)(MULT_SIZE-1) & MULT_16(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(71)<=signed(MULT_15(71)(MULT_SIZE-1) & MULT_15(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(71)(MULT_SIZE-1) & MULT_16(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(72)<=signed(MULT_15(72)(MULT_SIZE-1) & MULT_15(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(72)(MULT_SIZE-1) & MULT_16(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(73)<=signed(MULT_15(73)(MULT_SIZE-1) & MULT_15(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(73)(MULT_SIZE-1) & MULT_16(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(74)<=signed(MULT_15(74)(MULT_SIZE-1) & MULT_15(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(74)(MULT_SIZE-1) & MULT_16(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(75)<=signed(MULT_15(75)(MULT_SIZE-1) & MULT_15(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(75)(MULT_SIZE-1) & MULT_16(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(76)<=signed(MULT_15(76)(MULT_SIZE-1) & MULT_15(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(76)(MULT_SIZE-1) & MULT_16(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(77)<=signed(MULT_15(77)(MULT_SIZE-1) & MULT_15(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(77)(MULT_SIZE-1) & MULT_16(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(78)<=signed(MULT_15(78)(MULT_SIZE-1) & MULT_15(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(78)(MULT_SIZE-1) & MULT_16(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(79)<=signed(MULT_15(79)(MULT_SIZE-1) & MULT_15(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(79)(MULT_SIZE-1) & MULT_16(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(80)<=signed(MULT_15(80)(MULT_SIZE-1) & MULT_15(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(80)(MULT_SIZE-1) & MULT_16(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(81)<=signed(MULT_15(81)(MULT_SIZE-1) & MULT_15(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(81)(MULT_SIZE-1) & MULT_16(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(82)<=signed(MULT_15(82)(MULT_SIZE-1) & MULT_15(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(82)(MULT_SIZE-1) & MULT_16(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8(83)<=signed(MULT_15(83)(MULT_SIZE-1) & MULT_15(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_16(83)(MULT_SIZE-1) & MULT_16(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_9(0)<=signed(MULT_17(0)(MULT_SIZE-1) & MULT_17(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(0)(MULT_SIZE-1) & MULT_18(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(1)<=signed(MULT_17(1)(MULT_SIZE-1) & MULT_17(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(1)(MULT_SIZE-1) & MULT_18(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(2)<=signed(MULT_17(2)(MULT_SIZE-1) & MULT_17(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(2)(MULT_SIZE-1) & MULT_18(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(3)<=signed(MULT_17(3)(MULT_SIZE-1) & MULT_17(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(3)(MULT_SIZE-1) & MULT_18(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(4)<=signed(MULT_17(4)(MULT_SIZE-1) & MULT_17(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(4)(MULT_SIZE-1) & MULT_18(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(5)<=signed(MULT_17(5)(MULT_SIZE-1) & MULT_17(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(5)(MULT_SIZE-1) & MULT_18(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(6)<=signed(MULT_17(6)(MULT_SIZE-1) & MULT_17(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(6)(MULT_SIZE-1) & MULT_18(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(7)<=signed(MULT_17(7)(MULT_SIZE-1) & MULT_17(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(7)(MULT_SIZE-1) & MULT_18(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(8)<=signed(MULT_17(8)(MULT_SIZE-1) & MULT_17(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(8)(MULT_SIZE-1) & MULT_18(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(9)<=signed(MULT_17(9)(MULT_SIZE-1) & MULT_17(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(9)(MULT_SIZE-1) & MULT_18(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(10)<=signed(MULT_17(10)(MULT_SIZE-1) & MULT_17(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(10)(MULT_SIZE-1) & MULT_18(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(11)<=signed(MULT_17(11)(MULT_SIZE-1) & MULT_17(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(11)(MULT_SIZE-1) & MULT_18(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(12)<=signed(MULT_17(12)(MULT_SIZE-1) & MULT_17(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(12)(MULT_SIZE-1) & MULT_18(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(13)<=signed(MULT_17(13)(MULT_SIZE-1) & MULT_17(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(13)(MULT_SIZE-1) & MULT_18(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(14)<=signed(MULT_17(14)(MULT_SIZE-1) & MULT_17(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(14)(MULT_SIZE-1) & MULT_18(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(15)<=signed(MULT_17(15)(MULT_SIZE-1) & MULT_17(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(15)(MULT_SIZE-1) & MULT_18(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(16)<=signed(MULT_17(16)(MULT_SIZE-1) & MULT_17(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(16)(MULT_SIZE-1) & MULT_18(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(17)<=signed(MULT_17(17)(MULT_SIZE-1) & MULT_17(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(17)(MULT_SIZE-1) & MULT_18(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(18)<=signed(MULT_17(18)(MULT_SIZE-1) & MULT_17(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(18)(MULT_SIZE-1) & MULT_18(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(19)<=signed(MULT_17(19)(MULT_SIZE-1) & MULT_17(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(19)(MULT_SIZE-1) & MULT_18(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(20)<=signed(MULT_17(20)(MULT_SIZE-1) & MULT_17(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(20)(MULT_SIZE-1) & MULT_18(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(21)<=signed(MULT_17(21)(MULT_SIZE-1) & MULT_17(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(21)(MULT_SIZE-1) & MULT_18(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(22)<=signed(MULT_17(22)(MULT_SIZE-1) & MULT_17(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(22)(MULT_SIZE-1) & MULT_18(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(23)<=signed(MULT_17(23)(MULT_SIZE-1) & MULT_17(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(23)(MULT_SIZE-1) & MULT_18(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(24)<=signed(MULT_17(24)(MULT_SIZE-1) & MULT_17(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(24)(MULT_SIZE-1) & MULT_18(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(25)<=signed(MULT_17(25)(MULT_SIZE-1) & MULT_17(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(25)(MULT_SIZE-1) & MULT_18(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(26)<=signed(MULT_17(26)(MULT_SIZE-1) & MULT_17(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(26)(MULT_SIZE-1) & MULT_18(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(27)<=signed(MULT_17(27)(MULT_SIZE-1) & MULT_17(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(27)(MULT_SIZE-1) & MULT_18(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(28)<=signed(MULT_17(28)(MULT_SIZE-1) & MULT_17(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(28)(MULT_SIZE-1) & MULT_18(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(29)<=signed(MULT_17(29)(MULT_SIZE-1) & MULT_17(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(29)(MULT_SIZE-1) & MULT_18(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(30)<=signed(MULT_17(30)(MULT_SIZE-1) & MULT_17(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(30)(MULT_SIZE-1) & MULT_18(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(31)<=signed(MULT_17(31)(MULT_SIZE-1) & MULT_17(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(31)(MULT_SIZE-1) & MULT_18(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(32)<=signed(MULT_17(32)(MULT_SIZE-1) & MULT_17(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(32)(MULT_SIZE-1) & MULT_18(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(33)<=signed(MULT_17(33)(MULT_SIZE-1) & MULT_17(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(33)(MULT_SIZE-1) & MULT_18(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(34)<=signed(MULT_17(34)(MULT_SIZE-1) & MULT_17(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(34)(MULT_SIZE-1) & MULT_18(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(35)<=signed(MULT_17(35)(MULT_SIZE-1) & MULT_17(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(35)(MULT_SIZE-1) & MULT_18(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(36)<=signed(MULT_17(36)(MULT_SIZE-1) & MULT_17(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(36)(MULT_SIZE-1) & MULT_18(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(37)<=signed(MULT_17(37)(MULT_SIZE-1) & MULT_17(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(37)(MULT_SIZE-1) & MULT_18(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(38)<=signed(MULT_17(38)(MULT_SIZE-1) & MULT_17(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(38)(MULT_SIZE-1) & MULT_18(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(39)<=signed(MULT_17(39)(MULT_SIZE-1) & MULT_17(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(39)(MULT_SIZE-1) & MULT_18(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(40)<=signed(MULT_17(40)(MULT_SIZE-1) & MULT_17(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(40)(MULT_SIZE-1) & MULT_18(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(41)<=signed(MULT_17(41)(MULT_SIZE-1) & MULT_17(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(41)(MULT_SIZE-1) & MULT_18(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(42)<=signed(MULT_17(42)(MULT_SIZE-1) & MULT_17(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(42)(MULT_SIZE-1) & MULT_18(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(43)<=signed(MULT_17(43)(MULT_SIZE-1) & MULT_17(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(43)(MULT_SIZE-1) & MULT_18(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(44)<=signed(MULT_17(44)(MULT_SIZE-1) & MULT_17(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(44)(MULT_SIZE-1) & MULT_18(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(45)<=signed(MULT_17(45)(MULT_SIZE-1) & MULT_17(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(45)(MULT_SIZE-1) & MULT_18(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(46)<=signed(MULT_17(46)(MULT_SIZE-1) & MULT_17(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(46)(MULT_SIZE-1) & MULT_18(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(47)<=signed(MULT_17(47)(MULT_SIZE-1) & MULT_17(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(47)(MULT_SIZE-1) & MULT_18(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(48)<=signed(MULT_17(48)(MULT_SIZE-1) & MULT_17(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(48)(MULT_SIZE-1) & MULT_18(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(49)<=signed(MULT_17(49)(MULT_SIZE-1) & MULT_17(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(49)(MULT_SIZE-1) & MULT_18(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(50)<=signed(MULT_17(50)(MULT_SIZE-1) & MULT_17(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(50)(MULT_SIZE-1) & MULT_18(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(51)<=signed(MULT_17(51)(MULT_SIZE-1) & MULT_17(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(51)(MULT_SIZE-1) & MULT_18(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(52)<=signed(MULT_17(52)(MULT_SIZE-1) & MULT_17(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(52)(MULT_SIZE-1) & MULT_18(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(53)<=signed(MULT_17(53)(MULT_SIZE-1) & MULT_17(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(53)(MULT_SIZE-1) & MULT_18(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(54)<=signed(MULT_17(54)(MULT_SIZE-1) & MULT_17(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(54)(MULT_SIZE-1) & MULT_18(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(55)<=signed(MULT_17(55)(MULT_SIZE-1) & MULT_17(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(55)(MULT_SIZE-1) & MULT_18(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(56)<=signed(MULT_17(56)(MULT_SIZE-1) & MULT_17(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(56)(MULT_SIZE-1) & MULT_18(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(57)<=signed(MULT_17(57)(MULT_SIZE-1) & MULT_17(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(57)(MULT_SIZE-1) & MULT_18(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(58)<=signed(MULT_17(58)(MULT_SIZE-1) & MULT_17(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(58)(MULT_SIZE-1) & MULT_18(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(59)<=signed(MULT_17(59)(MULT_SIZE-1) & MULT_17(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(59)(MULT_SIZE-1) & MULT_18(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(60)<=signed(MULT_17(60)(MULT_SIZE-1) & MULT_17(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(60)(MULT_SIZE-1) & MULT_18(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(61)<=signed(MULT_17(61)(MULT_SIZE-1) & MULT_17(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(61)(MULT_SIZE-1) & MULT_18(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(62)<=signed(MULT_17(62)(MULT_SIZE-1) & MULT_17(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(62)(MULT_SIZE-1) & MULT_18(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(63)<=signed(MULT_17(63)(MULT_SIZE-1) & MULT_17(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(63)(MULT_SIZE-1) & MULT_18(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(64)<=signed(MULT_17(64)(MULT_SIZE-1) & MULT_17(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(64)(MULT_SIZE-1) & MULT_18(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(65)<=signed(MULT_17(65)(MULT_SIZE-1) & MULT_17(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(65)(MULT_SIZE-1) & MULT_18(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(66)<=signed(MULT_17(66)(MULT_SIZE-1) & MULT_17(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(66)(MULT_SIZE-1) & MULT_18(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(67)<=signed(MULT_17(67)(MULT_SIZE-1) & MULT_17(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(67)(MULT_SIZE-1) & MULT_18(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(68)<=signed(MULT_17(68)(MULT_SIZE-1) & MULT_17(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(68)(MULT_SIZE-1) & MULT_18(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(69)<=signed(MULT_17(69)(MULT_SIZE-1) & MULT_17(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(69)(MULT_SIZE-1) & MULT_18(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(70)<=signed(MULT_17(70)(MULT_SIZE-1) & MULT_17(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(70)(MULT_SIZE-1) & MULT_18(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(71)<=signed(MULT_17(71)(MULT_SIZE-1) & MULT_17(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(71)(MULT_SIZE-1) & MULT_18(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(72)<=signed(MULT_17(72)(MULT_SIZE-1) & MULT_17(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(72)(MULT_SIZE-1) & MULT_18(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(73)<=signed(MULT_17(73)(MULT_SIZE-1) & MULT_17(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(73)(MULT_SIZE-1) & MULT_18(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(74)<=signed(MULT_17(74)(MULT_SIZE-1) & MULT_17(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(74)(MULT_SIZE-1) & MULT_18(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(75)<=signed(MULT_17(75)(MULT_SIZE-1) & MULT_17(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(75)(MULT_SIZE-1) & MULT_18(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(76)<=signed(MULT_17(76)(MULT_SIZE-1) & MULT_17(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(76)(MULT_SIZE-1) & MULT_18(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(77)<=signed(MULT_17(77)(MULT_SIZE-1) & MULT_17(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(77)(MULT_SIZE-1) & MULT_18(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(78)<=signed(MULT_17(78)(MULT_SIZE-1) & MULT_17(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(78)(MULT_SIZE-1) & MULT_18(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(79)<=signed(MULT_17(79)(MULT_SIZE-1) & MULT_17(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(79)(MULT_SIZE-1) & MULT_18(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(80)<=signed(MULT_17(80)(MULT_SIZE-1) & MULT_17(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(80)(MULT_SIZE-1) & MULT_18(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(81)<=signed(MULT_17(81)(MULT_SIZE-1) & MULT_17(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(81)(MULT_SIZE-1) & MULT_18(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(82)<=signed(MULT_17(82)(MULT_SIZE-1) & MULT_17(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(82)(MULT_SIZE-1) & MULT_18(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9(83)<=signed(MULT_17(83)(MULT_SIZE-1) & MULT_17(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_18(83)(MULT_SIZE-1) & MULT_18(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_10(0)<=signed(MULT_19(0)(MULT_SIZE-1) & MULT_19(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(0)(MULT_SIZE-1) & MULT_20(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(1)<=signed(MULT_19(1)(MULT_SIZE-1) & MULT_19(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(1)(MULT_SIZE-1) & MULT_20(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(2)<=signed(MULT_19(2)(MULT_SIZE-1) & MULT_19(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(2)(MULT_SIZE-1) & MULT_20(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(3)<=signed(MULT_19(3)(MULT_SIZE-1) & MULT_19(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(3)(MULT_SIZE-1) & MULT_20(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(4)<=signed(MULT_19(4)(MULT_SIZE-1) & MULT_19(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(4)(MULT_SIZE-1) & MULT_20(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(5)<=signed(MULT_19(5)(MULT_SIZE-1) & MULT_19(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(5)(MULT_SIZE-1) & MULT_20(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(6)<=signed(MULT_19(6)(MULT_SIZE-1) & MULT_19(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(6)(MULT_SIZE-1) & MULT_20(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(7)<=signed(MULT_19(7)(MULT_SIZE-1) & MULT_19(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(7)(MULT_SIZE-1) & MULT_20(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(8)<=signed(MULT_19(8)(MULT_SIZE-1) & MULT_19(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(8)(MULT_SIZE-1) & MULT_20(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(9)<=signed(MULT_19(9)(MULT_SIZE-1) & MULT_19(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(9)(MULT_SIZE-1) & MULT_20(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(10)<=signed(MULT_19(10)(MULT_SIZE-1) & MULT_19(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(10)(MULT_SIZE-1) & MULT_20(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(11)<=signed(MULT_19(11)(MULT_SIZE-1) & MULT_19(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(11)(MULT_SIZE-1) & MULT_20(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(12)<=signed(MULT_19(12)(MULT_SIZE-1) & MULT_19(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(12)(MULT_SIZE-1) & MULT_20(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(13)<=signed(MULT_19(13)(MULT_SIZE-1) & MULT_19(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(13)(MULT_SIZE-1) & MULT_20(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(14)<=signed(MULT_19(14)(MULT_SIZE-1) & MULT_19(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(14)(MULT_SIZE-1) & MULT_20(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(15)<=signed(MULT_19(15)(MULT_SIZE-1) & MULT_19(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(15)(MULT_SIZE-1) & MULT_20(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(16)<=signed(MULT_19(16)(MULT_SIZE-1) & MULT_19(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(16)(MULT_SIZE-1) & MULT_20(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(17)<=signed(MULT_19(17)(MULT_SIZE-1) & MULT_19(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(17)(MULT_SIZE-1) & MULT_20(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(18)<=signed(MULT_19(18)(MULT_SIZE-1) & MULT_19(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(18)(MULT_SIZE-1) & MULT_20(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(19)<=signed(MULT_19(19)(MULT_SIZE-1) & MULT_19(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(19)(MULT_SIZE-1) & MULT_20(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(20)<=signed(MULT_19(20)(MULT_SIZE-1) & MULT_19(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(20)(MULT_SIZE-1) & MULT_20(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(21)<=signed(MULT_19(21)(MULT_SIZE-1) & MULT_19(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(21)(MULT_SIZE-1) & MULT_20(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(22)<=signed(MULT_19(22)(MULT_SIZE-1) & MULT_19(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(22)(MULT_SIZE-1) & MULT_20(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(23)<=signed(MULT_19(23)(MULT_SIZE-1) & MULT_19(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(23)(MULT_SIZE-1) & MULT_20(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(24)<=signed(MULT_19(24)(MULT_SIZE-1) & MULT_19(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(24)(MULT_SIZE-1) & MULT_20(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(25)<=signed(MULT_19(25)(MULT_SIZE-1) & MULT_19(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(25)(MULT_SIZE-1) & MULT_20(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(26)<=signed(MULT_19(26)(MULT_SIZE-1) & MULT_19(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(26)(MULT_SIZE-1) & MULT_20(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(27)<=signed(MULT_19(27)(MULT_SIZE-1) & MULT_19(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(27)(MULT_SIZE-1) & MULT_20(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(28)<=signed(MULT_19(28)(MULT_SIZE-1) & MULT_19(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(28)(MULT_SIZE-1) & MULT_20(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(29)<=signed(MULT_19(29)(MULT_SIZE-1) & MULT_19(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(29)(MULT_SIZE-1) & MULT_20(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(30)<=signed(MULT_19(30)(MULT_SIZE-1) & MULT_19(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(30)(MULT_SIZE-1) & MULT_20(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(31)<=signed(MULT_19(31)(MULT_SIZE-1) & MULT_19(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(31)(MULT_SIZE-1) & MULT_20(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(32)<=signed(MULT_19(32)(MULT_SIZE-1) & MULT_19(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(32)(MULT_SIZE-1) & MULT_20(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(33)<=signed(MULT_19(33)(MULT_SIZE-1) & MULT_19(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(33)(MULT_SIZE-1) & MULT_20(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(34)<=signed(MULT_19(34)(MULT_SIZE-1) & MULT_19(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(34)(MULT_SIZE-1) & MULT_20(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(35)<=signed(MULT_19(35)(MULT_SIZE-1) & MULT_19(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(35)(MULT_SIZE-1) & MULT_20(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(36)<=signed(MULT_19(36)(MULT_SIZE-1) & MULT_19(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(36)(MULT_SIZE-1) & MULT_20(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(37)<=signed(MULT_19(37)(MULT_SIZE-1) & MULT_19(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(37)(MULT_SIZE-1) & MULT_20(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(38)<=signed(MULT_19(38)(MULT_SIZE-1) & MULT_19(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(38)(MULT_SIZE-1) & MULT_20(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(39)<=signed(MULT_19(39)(MULT_SIZE-1) & MULT_19(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(39)(MULT_SIZE-1) & MULT_20(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(40)<=signed(MULT_19(40)(MULT_SIZE-1) & MULT_19(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(40)(MULT_SIZE-1) & MULT_20(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(41)<=signed(MULT_19(41)(MULT_SIZE-1) & MULT_19(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(41)(MULT_SIZE-1) & MULT_20(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(42)<=signed(MULT_19(42)(MULT_SIZE-1) & MULT_19(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(42)(MULT_SIZE-1) & MULT_20(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(43)<=signed(MULT_19(43)(MULT_SIZE-1) & MULT_19(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(43)(MULT_SIZE-1) & MULT_20(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(44)<=signed(MULT_19(44)(MULT_SIZE-1) & MULT_19(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(44)(MULT_SIZE-1) & MULT_20(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(45)<=signed(MULT_19(45)(MULT_SIZE-1) & MULT_19(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(45)(MULT_SIZE-1) & MULT_20(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(46)<=signed(MULT_19(46)(MULT_SIZE-1) & MULT_19(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(46)(MULT_SIZE-1) & MULT_20(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(47)<=signed(MULT_19(47)(MULT_SIZE-1) & MULT_19(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(47)(MULT_SIZE-1) & MULT_20(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(48)<=signed(MULT_19(48)(MULT_SIZE-1) & MULT_19(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(48)(MULT_SIZE-1) & MULT_20(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(49)<=signed(MULT_19(49)(MULT_SIZE-1) & MULT_19(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(49)(MULT_SIZE-1) & MULT_20(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(50)<=signed(MULT_19(50)(MULT_SIZE-1) & MULT_19(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(50)(MULT_SIZE-1) & MULT_20(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(51)<=signed(MULT_19(51)(MULT_SIZE-1) & MULT_19(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(51)(MULT_SIZE-1) & MULT_20(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(52)<=signed(MULT_19(52)(MULT_SIZE-1) & MULT_19(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(52)(MULT_SIZE-1) & MULT_20(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(53)<=signed(MULT_19(53)(MULT_SIZE-1) & MULT_19(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(53)(MULT_SIZE-1) & MULT_20(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(54)<=signed(MULT_19(54)(MULT_SIZE-1) & MULT_19(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(54)(MULT_SIZE-1) & MULT_20(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(55)<=signed(MULT_19(55)(MULT_SIZE-1) & MULT_19(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(55)(MULT_SIZE-1) & MULT_20(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(56)<=signed(MULT_19(56)(MULT_SIZE-1) & MULT_19(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(56)(MULT_SIZE-1) & MULT_20(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(57)<=signed(MULT_19(57)(MULT_SIZE-1) & MULT_19(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(57)(MULT_SIZE-1) & MULT_20(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(58)<=signed(MULT_19(58)(MULT_SIZE-1) & MULT_19(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(58)(MULT_SIZE-1) & MULT_20(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(59)<=signed(MULT_19(59)(MULT_SIZE-1) & MULT_19(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(59)(MULT_SIZE-1) & MULT_20(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(60)<=signed(MULT_19(60)(MULT_SIZE-1) & MULT_19(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(60)(MULT_SIZE-1) & MULT_20(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(61)<=signed(MULT_19(61)(MULT_SIZE-1) & MULT_19(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(61)(MULT_SIZE-1) & MULT_20(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(62)<=signed(MULT_19(62)(MULT_SIZE-1) & MULT_19(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(62)(MULT_SIZE-1) & MULT_20(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(63)<=signed(MULT_19(63)(MULT_SIZE-1) & MULT_19(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(63)(MULT_SIZE-1) & MULT_20(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(64)<=signed(MULT_19(64)(MULT_SIZE-1) & MULT_19(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(64)(MULT_SIZE-1) & MULT_20(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(65)<=signed(MULT_19(65)(MULT_SIZE-1) & MULT_19(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(65)(MULT_SIZE-1) & MULT_20(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(66)<=signed(MULT_19(66)(MULT_SIZE-1) & MULT_19(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(66)(MULT_SIZE-1) & MULT_20(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(67)<=signed(MULT_19(67)(MULT_SIZE-1) & MULT_19(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(67)(MULT_SIZE-1) & MULT_20(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(68)<=signed(MULT_19(68)(MULT_SIZE-1) & MULT_19(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(68)(MULT_SIZE-1) & MULT_20(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(69)<=signed(MULT_19(69)(MULT_SIZE-1) & MULT_19(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(69)(MULT_SIZE-1) & MULT_20(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(70)<=signed(MULT_19(70)(MULT_SIZE-1) & MULT_19(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(70)(MULT_SIZE-1) & MULT_20(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(71)<=signed(MULT_19(71)(MULT_SIZE-1) & MULT_19(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(71)(MULT_SIZE-1) & MULT_20(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(72)<=signed(MULT_19(72)(MULT_SIZE-1) & MULT_19(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(72)(MULT_SIZE-1) & MULT_20(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(73)<=signed(MULT_19(73)(MULT_SIZE-1) & MULT_19(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(73)(MULT_SIZE-1) & MULT_20(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(74)<=signed(MULT_19(74)(MULT_SIZE-1) & MULT_19(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(74)(MULT_SIZE-1) & MULT_20(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(75)<=signed(MULT_19(75)(MULT_SIZE-1) & MULT_19(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(75)(MULT_SIZE-1) & MULT_20(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(76)<=signed(MULT_19(76)(MULT_SIZE-1) & MULT_19(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(76)(MULT_SIZE-1) & MULT_20(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(77)<=signed(MULT_19(77)(MULT_SIZE-1) & MULT_19(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(77)(MULT_SIZE-1) & MULT_20(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(78)<=signed(MULT_19(78)(MULT_SIZE-1) & MULT_19(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(78)(MULT_SIZE-1) & MULT_20(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(79)<=signed(MULT_19(79)(MULT_SIZE-1) & MULT_19(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(79)(MULT_SIZE-1) & MULT_20(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(80)<=signed(MULT_19(80)(MULT_SIZE-1) & MULT_19(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(80)(MULT_SIZE-1) & MULT_20(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(81)<=signed(MULT_19(81)(MULT_SIZE-1) & MULT_19(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(81)(MULT_SIZE-1) & MULT_20(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(82)<=signed(MULT_19(82)(MULT_SIZE-1) & MULT_19(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(82)(MULT_SIZE-1) & MULT_20(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10(83)<=signed(MULT_19(83)(MULT_SIZE-1) & MULT_19(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_20(83)(MULT_SIZE-1) & MULT_20(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_11(0)<=signed(MULT_21(0)(MULT_SIZE-1) & MULT_21(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(0)(MULT_SIZE-1) & MULT_22(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(1)<=signed(MULT_21(1)(MULT_SIZE-1) & MULT_21(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(1)(MULT_SIZE-1) & MULT_22(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(2)<=signed(MULT_21(2)(MULT_SIZE-1) & MULT_21(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(2)(MULT_SIZE-1) & MULT_22(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(3)<=signed(MULT_21(3)(MULT_SIZE-1) & MULT_21(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(3)(MULT_SIZE-1) & MULT_22(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(4)<=signed(MULT_21(4)(MULT_SIZE-1) & MULT_21(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(4)(MULT_SIZE-1) & MULT_22(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(5)<=signed(MULT_21(5)(MULT_SIZE-1) & MULT_21(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(5)(MULT_SIZE-1) & MULT_22(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(6)<=signed(MULT_21(6)(MULT_SIZE-1) & MULT_21(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(6)(MULT_SIZE-1) & MULT_22(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(7)<=signed(MULT_21(7)(MULT_SIZE-1) & MULT_21(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(7)(MULT_SIZE-1) & MULT_22(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(8)<=signed(MULT_21(8)(MULT_SIZE-1) & MULT_21(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(8)(MULT_SIZE-1) & MULT_22(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(9)<=signed(MULT_21(9)(MULT_SIZE-1) & MULT_21(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(9)(MULT_SIZE-1) & MULT_22(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(10)<=signed(MULT_21(10)(MULT_SIZE-1) & MULT_21(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(10)(MULT_SIZE-1) & MULT_22(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(11)<=signed(MULT_21(11)(MULT_SIZE-1) & MULT_21(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(11)(MULT_SIZE-1) & MULT_22(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(12)<=signed(MULT_21(12)(MULT_SIZE-1) & MULT_21(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(12)(MULT_SIZE-1) & MULT_22(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(13)<=signed(MULT_21(13)(MULT_SIZE-1) & MULT_21(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(13)(MULT_SIZE-1) & MULT_22(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(14)<=signed(MULT_21(14)(MULT_SIZE-1) & MULT_21(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(14)(MULT_SIZE-1) & MULT_22(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(15)<=signed(MULT_21(15)(MULT_SIZE-1) & MULT_21(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(15)(MULT_SIZE-1) & MULT_22(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(16)<=signed(MULT_21(16)(MULT_SIZE-1) & MULT_21(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(16)(MULT_SIZE-1) & MULT_22(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(17)<=signed(MULT_21(17)(MULT_SIZE-1) & MULT_21(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(17)(MULT_SIZE-1) & MULT_22(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(18)<=signed(MULT_21(18)(MULT_SIZE-1) & MULT_21(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(18)(MULT_SIZE-1) & MULT_22(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(19)<=signed(MULT_21(19)(MULT_SIZE-1) & MULT_21(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(19)(MULT_SIZE-1) & MULT_22(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(20)<=signed(MULT_21(20)(MULT_SIZE-1) & MULT_21(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(20)(MULT_SIZE-1) & MULT_22(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(21)<=signed(MULT_21(21)(MULT_SIZE-1) & MULT_21(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(21)(MULT_SIZE-1) & MULT_22(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(22)<=signed(MULT_21(22)(MULT_SIZE-1) & MULT_21(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(22)(MULT_SIZE-1) & MULT_22(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(23)<=signed(MULT_21(23)(MULT_SIZE-1) & MULT_21(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(23)(MULT_SIZE-1) & MULT_22(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(24)<=signed(MULT_21(24)(MULT_SIZE-1) & MULT_21(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(24)(MULT_SIZE-1) & MULT_22(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(25)<=signed(MULT_21(25)(MULT_SIZE-1) & MULT_21(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(25)(MULT_SIZE-1) & MULT_22(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(26)<=signed(MULT_21(26)(MULT_SIZE-1) & MULT_21(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(26)(MULT_SIZE-1) & MULT_22(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(27)<=signed(MULT_21(27)(MULT_SIZE-1) & MULT_21(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(27)(MULT_SIZE-1) & MULT_22(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(28)<=signed(MULT_21(28)(MULT_SIZE-1) & MULT_21(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(28)(MULT_SIZE-1) & MULT_22(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(29)<=signed(MULT_21(29)(MULT_SIZE-1) & MULT_21(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(29)(MULT_SIZE-1) & MULT_22(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(30)<=signed(MULT_21(30)(MULT_SIZE-1) & MULT_21(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(30)(MULT_SIZE-1) & MULT_22(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(31)<=signed(MULT_21(31)(MULT_SIZE-1) & MULT_21(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(31)(MULT_SIZE-1) & MULT_22(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(32)<=signed(MULT_21(32)(MULT_SIZE-1) & MULT_21(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(32)(MULT_SIZE-1) & MULT_22(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(33)<=signed(MULT_21(33)(MULT_SIZE-1) & MULT_21(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(33)(MULT_SIZE-1) & MULT_22(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(34)<=signed(MULT_21(34)(MULT_SIZE-1) & MULT_21(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(34)(MULT_SIZE-1) & MULT_22(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(35)<=signed(MULT_21(35)(MULT_SIZE-1) & MULT_21(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(35)(MULT_SIZE-1) & MULT_22(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(36)<=signed(MULT_21(36)(MULT_SIZE-1) & MULT_21(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(36)(MULT_SIZE-1) & MULT_22(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(37)<=signed(MULT_21(37)(MULT_SIZE-1) & MULT_21(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(37)(MULT_SIZE-1) & MULT_22(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(38)<=signed(MULT_21(38)(MULT_SIZE-1) & MULT_21(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(38)(MULT_SIZE-1) & MULT_22(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(39)<=signed(MULT_21(39)(MULT_SIZE-1) & MULT_21(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(39)(MULT_SIZE-1) & MULT_22(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(40)<=signed(MULT_21(40)(MULT_SIZE-1) & MULT_21(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(40)(MULT_SIZE-1) & MULT_22(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(41)<=signed(MULT_21(41)(MULT_SIZE-1) & MULT_21(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(41)(MULT_SIZE-1) & MULT_22(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(42)<=signed(MULT_21(42)(MULT_SIZE-1) & MULT_21(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(42)(MULT_SIZE-1) & MULT_22(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(43)<=signed(MULT_21(43)(MULT_SIZE-1) & MULT_21(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(43)(MULT_SIZE-1) & MULT_22(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(44)<=signed(MULT_21(44)(MULT_SIZE-1) & MULT_21(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(44)(MULT_SIZE-1) & MULT_22(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(45)<=signed(MULT_21(45)(MULT_SIZE-1) & MULT_21(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(45)(MULT_SIZE-1) & MULT_22(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(46)<=signed(MULT_21(46)(MULT_SIZE-1) & MULT_21(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(46)(MULT_SIZE-1) & MULT_22(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(47)<=signed(MULT_21(47)(MULT_SIZE-1) & MULT_21(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(47)(MULT_SIZE-1) & MULT_22(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(48)<=signed(MULT_21(48)(MULT_SIZE-1) & MULT_21(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(48)(MULT_SIZE-1) & MULT_22(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(49)<=signed(MULT_21(49)(MULT_SIZE-1) & MULT_21(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(49)(MULT_SIZE-1) & MULT_22(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(50)<=signed(MULT_21(50)(MULT_SIZE-1) & MULT_21(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(50)(MULT_SIZE-1) & MULT_22(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(51)<=signed(MULT_21(51)(MULT_SIZE-1) & MULT_21(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(51)(MULT_SIZE-1) & MULT_22(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(52)<=signed(MULT_21(52)(MULT_SIZE-1) & MULT_21(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(52)(MULT_SIZE-1) & MULT_22(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(53)<=signed(MULT_21(53)(MULT_SIZE-1) & MULT_21(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(53)(MULT_SIZE-1) & MULT_22(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(54)<=signed(MULT_21(54)(MULT_SIZE-1) & MULT_21(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(54)(MULT_SIZE-1) & MULT_22(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(55)<=signed(MULT_21(55)(MULT_SIZE-1) & MULT_21(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(55)(MULT_SIZE-1) & MULT_22(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(56)<=signed(MULT_21(56)(MULT_SIZE-1) & MULT_21(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(56)(MULT_SIZE-1) & MULT_22(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(57)<=signed(MULT_21(57)(MULT_SIZE-1) & MULT_21(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(57)(MULT_SIZE-1) & MULT_22(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(58)<=signed(MULT_21(58)(MULT_SIZE-1) & MULT_21(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(58)(MULT_SIZE-1) & MULT_22(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(59)<=signed(MULT_21(59)(MULT_SIZE-1) & MULT_21(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(59)(MULT_SIZE-1) & MULT_22(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(60)<=signed(MULT_21(60)(MULT_SIZE-1) & MULT_21(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(60)(MULT_SIZE-1) & MULT_22(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(61)<=signed(MULT_21(61)(MULT_SIZE-1) & MULT_21(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(61)(MULT_SIZE-1) & MULT_22(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(62)<=signed(MULT_21(62)(MULT_SIZE-1) & MULT_21(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(62)(MULT_SIZE-1) & MULT_22(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(63)<=signed(MULT_21(63)(MULT_SIZE-1) & MULT_21(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(63)(MULT_SIZE-1) & MULT_22(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(64)<=signed(MULT_21(64)(MULT_SIZE-1) & MULT_21(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(64)(MULT_SIZE-1) & MULT_22(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(65)<=signed(MULT_21(65)(MULT_SIZE-1) & MULT_21(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(65)(MULT_SIZE-1) & MULT_22(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(66)<=signed(MULT_21(66)(MULT_SIZE-1) & MULT_21(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(66)(MULT_SIZE-1) & MULT_22(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(67)<=signed(MULT_21(67)(MULT_SIZE-1) & MULT_21(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(67)(MULT_SIZE-1) & MULT_22(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(68)<=signed(MULT_21(68)(MULT_SIZE-1) & MULT_21(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(68)(MULT_SIZE-1) & MULT_22(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(69)<=signed(MULT_21(69)(MULT_SIZE-1) & MULT_21(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(69)(MULT_SIZE-1) & MULT_22(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(70)<=signed(MULT_21(70)(MULT_SIZE-1) & MULT_21(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(70)(MULT_SIZE-1) & MULT_22(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(71)<=signed(MULT_21(71)(MULT_SIZE-1) & MULT_21(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(71)(MULT_SIZE-1) & MULT_22(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(72)<=signed(MULT_21(72)(MULT_SIZE-1) & MULT_21(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(72)(MULT_SIZE-1) & MULT_22(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(73)<=signed(MULT_21(73)(MULT_SIZE-1) & MULT_21(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(73)(MULT_SIZE-1) & MULT_22(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(74)<=signed(MULT_21(74)(MULT_SIZE-1) & MULT_21(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(74)(MULT_SIZE-1) & MULT_22(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(75)<=signed(MULT_21(75)(MULT_SIZE-1) & MULT_21(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(75)(MULT_SIZE-1) & MULT_22(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(76)<=signed(MULT_21(76)(MULT_SIZE-1) & MULT_21(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(76)(MULT_SIZE-1) & MULT_22(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(77)<=signed(MULT_21(77)(MULT_SIZE-1) & MULT_21(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(77)(MULT_SIZE-1) & MULT_22(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(78)<=signed(MULT_21(78)(MULT_SIZE-1) & MULT_21(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(78)(MULT_SIZE-1) & MULT_22(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(79)<=signed(MULT_21(79)(MULT_SIZE-1) & MULT_21(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(79)(MULT_SIZE-1) & MULT_22(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(80)<=signed(MULT_21(80)(MULT_SIZE-1) & MULT_21(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(80)(MULT_SIZE-1) & MULT_22(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(81)<=signed(MULT_21(81)(MULT_SIZE-1) & MULT_21(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(81)(MULT_SIZE-1) & MULT_22(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(82)<=signed(MULT_21(82)(MULT_SIZE-1) & MULT_21(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(82)(MULT_SIZE-1) & MULT_22(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11(83)<=signed(MULT_21(83)(MULT_SIZE-1) & MULT_21(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_22(83)(MULT_SIZE-1) & MULT_22(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_12(0)<=signed(MULT_23(0)(MULT_SIZE-1) & MULT_23(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(0)(MULT_SIZE-1) & MULT_24(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(1)<=signed(MULT_23(1)(MULT_SIZE-1) & MULT_23(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(1)(MULT_SIZE-1) & MULT_24(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(2)<=signed(MULT_23(2)(MULT_SIZE-1) & MULT_23(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(2)(MULT_SIZE-1) & MULT_24(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(3)<=signed(MULT_23(3)(MULT_SIZE-1) & MULT_23(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(3)(MULT_SIZE-1) & MULT_24(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(4)<=signed(MULT_23(4)(MULT_SIZE-1) & MULT_23(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(4)(MULT_SIZE-1) & MULT_24(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(5)<=signed(MULT_23(5)(MULT_SIZE-1) & MULT_23(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(5)(MULT_SIZE-1) & MULT_24(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(6)<=signed(MULT_23(6)(MULT_SIZE-1) & MULT_23(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(6)(MULT_SIZE-1) & MULT_24(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(7)<=signed(MULT_23(7)(MULT_SIZE-1) & MULT_23(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(7)(MULT_SIZE-1) & MULT_24(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(8)<=signed(MULT_23(8)(MULT_SIZE-1) & MULT_23(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(8)(MULT_SIZE-1) & MULT_24(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(9)<=signed(MULT_23(9)(MULT_SIZE-1) & MULT_23(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(9)(MULT_SIZE-1) & MULT_24(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(10)<=signed(MULT_23(10)(MULT_SIZE-1) & MULT_23(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(10)(MULT_SIZE-1) & MULT_24(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(11)<=signed(MULT_23(11)(MULT_SIZE-1) & MULT_23(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(11)(MULT_SIZE-1) & MULT_24(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(12)<=signed(MULT_23(12)(MULT_SIZE-1) & MULT_23(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(12)(MULT_SIZE-1) & MULT_24(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(13)<=signed(MULT_23(13)(MULT_SIZE-1) & MULT_23(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(13)(MULT_SIZE-1) & MULT_24(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(14)<=signed(MULT_23(14)(MULT_SIZE-1) & MULT_23(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(14)(MULT_SIZE-1) & MULT_24(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(15)<=signed(MULT_23(15)(MULT_SIZE-1) & MULT_23(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(15)(MULT_SIZE-1) & MULT_24(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(16)<=signed(MULT_23(16)(MULT_SIZE-1) & MULT_23(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(16)(MULT_SIZE-1) & MULT_24(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(17)<=signed(MULT_23(17)(MULT_SIZE-1) & MULT_23(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(17)(MULT_SIZE-1) & MULT_24(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(18)<=signed(MULT_23(18)(MULT_SIZE-1) & MULT_23(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(18)(MULT_SIZE-1) & MULT_24(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(19)<=signed(MULT_23(19)(MULT_SIZE-1) & MULT_23(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(19)(MULT_SIZE-1) & MULT_24(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(20)<=signed(MULT_23(20)(MULT_SIZE-1) & MULT_23(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(20)(MULT_SIZE-1) & MULT_24(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(21)<=signed(MULT_23(21)(MULT_SIZE-1) & MULT_23(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(21)(MULT_SIZE-1) & MULT_24(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(22)<=signed(MULT_23(22)(MULT_SIZE-1) & MULT_23(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(22)(MULT_SIZE-1) & MULT_24(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(23)<=signed(MULT_23(23)(MULT_SIZE-1) & MULT_23(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(23)(MULT_SIZE-1) & MULT_24(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(24)<=signed(MULT_23(24)(MULT_SIZE-1) & MULT_23(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(24)(MULT_SIZE-1) & MULT_24(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(25)<=signed(MULT_23(25)(MULT_SIZE-1) & MULT_23(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(25)(MULT_SIZE-1) & MULT_24(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(26)<=signed(MULT_23(26)(MULT_SIZE-1) & MULT_23(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(26)(MULT_SIZE-1) & MULT_24(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(27)<=signed(MULT_23(27)(MULT_SIZE-1) & MULT_23(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(27)(MULT_SIZE-1) & MULT_24(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(28)<=signed(MULT_23(28)(MULT_SIZE-1) & MULT_23(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(28)(MULT_SIZE-1) & MULT_24(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(29)<=signed(MULT_23(29)(MULT_SIZE-1) & MULT_23(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(29)(MULT_SIZE-1) & MULT_24(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(30)<=signed(MULT_23(30)(MULT_SIZE-1) & MULT_23(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(30)(MULT_SIZE-1) & MULT_24(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(31)<=signed(MULT_23(31)(MULT_SIZE-1) & MULT_23(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(31)(MULT_SIZE-1) & MULT_24(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(32)<=signed(MULT_23(32)(MULT_SIZE-1) & MULT_23(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(32)(MULT_SIZE-1) & MULT_24(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(33)<=signed(MULT_23(33)(MULT_SIZE-1) & MULT_23(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(33)(MULT_SIZE-1) & MULT_24(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(34)<=signed(MULT_23(34)(MULT_SIZE-1) & MULT_23(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(34)(MULT_SIZE-1) & MULT_24(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(35)<=signed(MULT_23(35)(MULT_SIZE-1) & MULT_23(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(35)(MULT_SIZE-1) & MULT_24(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(36)<=signed(MULT_23(36)(MULT_SIZE-1) & MULT_23(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(36)(MULT_SIZE-1) & MULT_24(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(37)<=signed(MULT_23(37)(MULT_SIZE-1) & MULT_23(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(37)(MULT_SIZE-1) & MULT_24(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(38)<=signed(MULT_23(38)(MULT_SIZE-1) & MULT_23(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(38)(MULT_SIZE-1) & MULT_24(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(39)<=signed(MULT_23(39)(MULT_SIZE-1) & MULT_23(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(39)(MULT_SIZE-1) & MULT_24(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(40)<=signed(MULT_23(40)(MULT_SIZE-1) & MULT_23(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(40)(MULT_SIZE-1) & MULT_24(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(41)<=signed(MULT_23(41)(MULT_SIZE-1) & MULT_23(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(41)(MULT_SIZE-1) & MULT_24(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(42)<=signed(MULT_23(42)(MULT_SIZE-1) & MULT_23(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(42)(MULT_SIZE-1) & MULT_24(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(43)<=signed(MULT_23(43)(MULT_SIZE-1) & MULT_23(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(43)(MULT_SIZE-1) & MULT_24(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(44)<=signed(MULT_23(44)(MULT_SIZE-1) & MULT_23(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(44)(MULT_SIZE-1) & MULT_24(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(45)<=signed(MULT_23(45)(MULT_SIZE-1) & MULT_23(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(45)(MULT_SIZE-1) & MULT_24(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(46)<=signed(MULT_23(46)(MULT_SIZE-1) & MULT_23(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(46)(MULT_SIZE-1) & MULT_24(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(47)<=signed(MULT_23(47)(MULT_SIZE-1) & MULT_23(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(47)(MULT_SIZE-1) & MULT_24(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(48)<=signed(MULT_23(48)(MULT_SIZE-1) & MULT_23(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(48)(MULT_SIZE-1) & MULT_24(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(49)<=signed(MULT_23(49)(MULT_SIZE-1) & MULT_23(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(49)(MULT_SIZE-1) & MULT_24(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(50)<=signed(MULT_23(50)(MULT_SIZE-1) & MULT_23(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(50)(MULT_SIZE-1) & MULT_24(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(51)<=signed(MULT_23(51)(MULT_SIZE-1) & MULT_23(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(51)(MULT_SIZE-1) & MULT_24(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(52)<=signed(MULT_23(52)(MULT_SIZE-1) & MULT_23(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(52)(MULT_SIZE-1) & MULT_24(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(53)<=signed(MULT_23(53)(MULT_SIZE-1) & MULT_23(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(53)(MULT_SIZE-1) & MULT_24(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(54)<=signed(MULT_23(54)(MULT_SIZE-1) & MULT_23(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(54)(MULT_SIZE-1) & MULT_24(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(55)<=signed(MULT_23(55)(MULT_SIZE-1) & MULT_23(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(55)(MULT_SIZE-1) & MULT_24(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(56)<=signed(MULT_23(56)(MULT_SIZE-1) & MULT_23(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(56)(MULT_SIZE-1) & MULT_24(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(57)<=signed(MULT_23(57)(MULT_SIZE-1) & MULT_23(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(57)(MULT_SIZE-1) & MULT_24(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(58)<=signed(MULT_23(58)(MULT_SIZE-1) & MULT_23(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(58)(MULT_SIZE-1) & MULT_24(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(59)<=signed(MULT_23(59)(MULT_SIZE-1) & MULT_23(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(59)(MULT_SIZE-1) & MULT_24(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(60)<=signed(MULT_23(60)(MULT_SIZE-1) & MULT_23(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(60)(MULT_SIZE-1) & MULT_24(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(61)<=signed(MULT_23(61)(MULT_SIZE-1) & MULT_23(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(61)(MULT_SIZE-1) & MULT_24(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(62)<=signed(MULT_23(62)(MULT_SIZE-1) & MULT_23(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(62)(MULT_SIZE-1) & MULT_24(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(63)<=signed(MULT_23(63)(MULT_SIZE-1) & MULT_23(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(63)(MULT_SIZE-1) & MULT_24(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(64)<=signed(MULT_23(64)(MULT_SIZE-1) & MULT_23(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(64)(MULT_SIZE-1) & MULT_24(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(65)<=signed(MULT_23(65)(MULT_SIZE-1) & MULT_23(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(65)(MULT_SIZE-1) & MULT_24(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(66)<=signed(MULT_23(66)(MULT_SIZE-1) & MULT_23(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(66)(MULT_SIZE-1) & MULT_24(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(67)<=signed(MULT_23(67)(MULT_SIZE-1) & MULT_23(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(67)(MULT_SIZE-1) & MULT_24(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(68)<=signed(MULT_23(68)(MULT_SIZE-1) & MULT_23(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(68)(MULT_SIZE-1) & MULT_24(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(69)<=signed(MULT_23(69)(MULT_SIZE-1) & MULT_23(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(69)(MULT_SIZE-1) & MULT_24(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(70)<=signed(MULT_23(70)(MULT_SIZE-1) & MULT_23(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(70)(MULT_SIZE-1) & MULT_24(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(71)<=signed(MULT_23(71)(MULT_SIZE-1) & MULT_23(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(71)(MULT_SIZE-1) & MULT_24(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(72)<=signed(MULT_23(72)(MULT_SIZE-1) & MULT_23(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(72)(MULT_SIZE-1) & MULT_24(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(73)<=signed(MULT_23(73)(MULT_SIZE-1) & MULT_23(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(73)(MULT_SIZE-1) & MULT_24(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(74)<=signed(MULT_23(74)(MULT_SIZE-1) & MULT_23(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(74)(MULT_SIZE-1) & MULT_24(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(75)<=signed(MULT_23(75)(MULT_SIZE-1) & MULT_23(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(75)(MULT_SIZE-1) & MULT_24(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(76)<=signed(MULT_23(76)(MULT_SIZE-1) & MULT_23(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(76)(MULT_SIZE-1) & MULT_24(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(77)<=signed(MULT_23(77)(MULT_SIZE-1) & MULT_23(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(77)(MULT_SIZE-1) & MULT_24(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(78)<=signed(MULT_23(78)(MULT_SIZE-1) & MULT_23(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(78)(MULT_SIZE-1) & MULT_24(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(79)<=signed(MULT_23(79)(MULT_SIZE-1) & MULT_23(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(79)(MULT_SIZE-1) & MULT_24(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(80)<=signed(MULT_23(80)(MULT_SIZE-1) & MULT_23(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(80)(MULT_SIZE-1) & MULT_24(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(81)<=signed(MULT_23(81)(MULT_SIZE-1) & MULT_23(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(81)(MULT_SIZE-1) & MULT_24(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(82)<=signed(MULT_23(82)(MULT_SIZE-1) & MULT_23(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(82)(MULT_SIZE-1) & MULT_24(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12(83)<=signed(MULT_23(83)(MULT_SIZE-1) & MULT_23(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_24(83)(MULT_SIZE-1) & MULT_24(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_13(0)<=signed(MULT_25(0)(MULT_SIZE-1) & MULT_25(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(0)(MULT_SIZE-1) & MULT_26(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(1)<=signed(MULT_25(1)(MULT_SIZE-1) & MULT_25(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(1)(MULT_SIZE-1) & MULT_26(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(2)<=signed(MULT_25(2)(MULT_SIZE-1) & MULT_25(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(2)(MULT_SIZE-1) & MULT_26(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(3)<=signed(MULT_25(3)(MULT_SIZE-1) & MULT_25(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(3)(MULT_SIZE-1) & MULT_26(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(4)<=signed(MULT_25(4)(MULT_SIZE-1) & MULT_25(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(4)(MULT_SIZE-1) & MULT_26(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(5)<=signed(MULT_25(5)(MULT_SIZE-1) & MULT_25(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(5)(MULT_SIZE-1) & MULT_26(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(6)<=signed(MULT_25(6)(MULT_SIZE-1) & MULT_25(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(6)(MULT_SIZE-1) & MULT_26(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(7)<=signed(MULT_25(7)(MULT_SIZE-1) & MULT_25(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(7)(MULT_SIZE-1) & MULT_26(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(8)<=signed(MULT_25(8)(MULT_SIZE-1) & MULT_25(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(8)(MULT_SIZE-1) & MULT_26(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(9)<=signed(MULT_25(9)(MULT_SIZE-1) & MULT_25(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(9)(MULT_SIZE-1) & MULT_26(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(10)<=signed(MULT_25(10)(MULT_SIZE-1) & MULT_25(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(10)(MULT_SIZE-1) & MULT_26(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(11)<=signed(MULT_25(11)(MULT_SIZE-1) & MULT_25(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(11)(MULT_SIZE-1) & MULT_26(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(12)<=signed(MULT_25(12)(MULT_SIZE-1) & MULT_25(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(12)(MULT_SIZE-1) & MULT_26(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(13)<=signed(MULT_25(13)(MULT_SIZE-1) & MULT_25(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(13)(MULT_SIZE-1) & MULT_26(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(14)<=signed(MULT_25(14)(MULT_SIZE-1) & MULT_25(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(14)(MULT_SIZE-1) & MULT_26(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(15)<=signed(MULT_25(15)(MULT_SIZE-1) & MULT_25(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(15)(MULT_SIZE-1) & MULT_26(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(16)<=signed(MULT_25(16)(MULT_SIZE-1) & MULT_25(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(16)(MULT_SIZE-1) & MULT_26(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(17)<=signed(MULT_25(17)(MULT_SIZE-1) & MULT_25(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(17)(MULT_SIZE-1) & MULT_26(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(18)<=signed(MULT_25(18)(MULT_SIZE-1) & MULT_25(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(18)(MULT_SIZE-1) & MULT_26(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(19)<=signed(MULT_25(19)(MULT_SIZE-1) & MULT_25(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(19)(MULT_SIZE-1) & MULT_26(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(20)<=signed(MULT_25(20)(MULT_SIZE-1) & MULT_25(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(20)(MULT_SIZE-1) & MULT_26(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(21)<=signed(MULT_25(21)(MULT_SIZE-1) & MULT_25(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(21)(MULT_SIZE-1) & MULT_26(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(22)<=signed(MULT_25(22)(MULT_SIZE-1) & MULT_25(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(22)(MULT_SIZE-1) & MULT_26(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(23)<=signed(MULT_25(23)(MULT_SIZE-1) & MULT_25(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(23)(MULT_SIZE-1) & MULT_26(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(24)<=signed(MULT_25(24)(MULT_SIZE-1) & MULT_25(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(24)(MULT_SIZE-1) & MULT_26(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(25)<=signed(MULT_25(25)(MULT_SIZE-1) & MULT_25(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(25)(MULT_SIZE-1) & MULT_26(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(26)<=signed(MULT_25(26)(MULT_SIZE-1) & MULT_25(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(26)(MULT_SIZE-1) & MULT_26(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(27)<=signed(MULT_25(27)(MULT_SIZE-1) & MULT_25(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(27)(MULT_SIZE-1) & MULT_26(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(28)<=signed(MULT_25(28)(MULT_SIZE-1) & MULT_25(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(28)(MULT_SIZE-1) & MULT_26(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(29)<=signed(MULT_25(29)(MULT_SIZE-1) & MULT_25(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(29)(MULT_SIZE-1) & MULT_26(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(30)<=signed(MULT_25(30)(MULT_SIZE-1) & MULT_25(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(30)(MULT_SIZE-1) & MULT_26(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(31)<=signed(MULT_25(31)(MULT_SIZE-1) & MULT_25(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(31)(MULT_SIZE-1) & MULT_26(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(32)<=signed(MULT_25(32)(MULT_SIZE-1) & MULT_25(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(32)(MULT_SIZE-1) & MULT_26(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(33)<=signed(MULT_25(33)(MULT_SIZE-1) & MULT_25(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(33)(MULT_SIZE-1) & MULT_26(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(34)<=signed(MULT_25(34)(MULT_SIZE-1) & MULT_25(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(34)(MULT_SIZE-1) & MULT_26(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(35)<=signed(MULT_25(35)(MULT_SIZE-1) & MULT_25(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(35)(MULT_SIZE-1) & MULT_26(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(36)<=signed(MULT_25(36)(MULT_SIZE-1) & MULT_25(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(36)(MULT_SIZE-1) & MULT_26(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(37)<=signed(MULT_25(37)(MULT_SIZE-1) & MULT_25(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(37)(MULT_SIZE-1) & MULT_26(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(38)<=signed(MULT_25(38)(MULT_SIZE-1) & MULT_25(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(38)(MULT_SIZE-1) & MULT_26(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(39)<=signed(MULT_25(39)(MULT_SIZE-1) & MULT_25(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(39)(MULT_SIZE-1) & MULT_26(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(40)<=signed(MULT_25(40)(MULT_SIZE-1) & MULT_25(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(40)(MULT_SIZE-1) & MULT_26(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(41)<=signed(MULT_25(41)(MULT_SIZE-1) & MULT_25(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(41)(MULT_SIZE-1) & MULT_26(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(42)<=signed(MULT_25(42)(MULT_SIZE-1) & MULT_25(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(42)(MULT_SIZE-1) & MULT_26(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(43)<=signed(MULT_25(43)(MULT_SIZE-1) & MULT_25(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(43)(MULT_SIZE-1) & MULT_26(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(44)<=signed(MULT_25(44)(MULT_SIZE-1) & MULT_25(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(44)(MULT_SIZE-1) & MULT_26(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(45)<=signed(MULT_25(45)(MULT_SIZE-1) & MULT_25(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(45)(MULT_SIZE-1) & MULT_26(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(46)<=signed(MULT_25(46)(MULT_SIZE-1) & MULT_25(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(46)(MULT_SIZE-1) & MULT_26(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(47)<=signed(MULT_25(47)(MULT_SIZE-1) & MULT_25(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(47)(MULT_SIZE-1) & MULT_26(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(48)<=signed(MULT_25(48)(MULT_SIZE-1) & MULT_25(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(48)(MULT_SIZE-1) & MULT_26(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(49)<=signed(MULT_25(49)(MULT_SIZE-1) & MULT_25(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(49)(MULT_SIZE-1) & MULT_26(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(50)<=signed(MULT_25(50)(MULT_SIZE-1) & MULT_25(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(50)(MULT_SIZE-1) & MULT_26(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(51)<=signed(MULT_25(51)(MULT_SIZE-1) & MULT_25(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(51)(MULT_SIZE-1) & MULT_26(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(52)<=signed(MULT_25(52)(MULT_SIZE-1) & MULT_25(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(52)(MULT_SIZE-1) & MULT_26(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(53)<=signed(MULT_25(53)(MULT_SIZE-1) & MULT_25(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(53)(MULT_SIZE-1) & MULT_26(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(54)<=signed(MULT_25(54)(MULT_SIZE-1) & MULT_25(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(54)(MULT_SIZE-1) & MULT_26(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(55)<=signed(MULT_25(55)(MULT_SIZE-1) & MULT_25(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(55)(MULT_SIZE-1) & MULT_26(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(56)<=signed(MULT_25(56)(MULT_SIZE-1) & MULT_25(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(56)(MULT_SIZE-1) & MULT_26(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(57)<=signed(MULT_25(57)(MULT_SIZE-1) & MULT_25(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(57)(MULT_SIZE-1) & MULT_26(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(58)<=signed(MULT_25(58)(MULT_SIZE-1) & MULT_25(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(58)(MULT_SIZE-1) & MULT_26(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(59)<=signed(MULT_25(59)(MULT_SIZE-1) & MULT_25(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(59)(MULT_SIZE-1) & MULT_26(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(60)<=signed(MULT_25(60)(MULT_SIZE-1) & MULT_25(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(60)(MULT_SIZE-1) & MULT_26(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(61)<=signed(MULT_25(61)(MULT_SIZE-1) & MULT_25(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(61)(MULT_SIZE-1) & MULT_26(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(62)<=signed(MULT_25(62)(MULT_SIZE-1) & MULT_25(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(62)(MULT_SIZE-1) & MULT_26(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(63)<=signed(MULT_25(63)(MULT_SIZE-1) & MULT_25(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(63)(MULT_SIZE-1) & MULT_26(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(64)<=signed(MULT_25(64)(MULT_SIZE-1) & MULT_25(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(64)(MULT_SIZE-1) & MULT_26(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(65)<=signed(MULT_25(65)(MULT_SIZE-1) & MULT_25(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(65)(MULT_SIZE-1) & MULT_26(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(66)<=signed(MULT_25(66)(MULT_SIZE-1) & MULT_25(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(66)(MULT_SIZE-1) & MULT_26(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(67)<=signed(MULT_25(67)(MULT_SIZE-1) & MULT_25(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(67)(MULT_SIZE-1) & MULT_26(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(68)<=signed(MULT_25(68)(MULT_SIZE-1) & MULT_25(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(68)(MULT_SIZE-1) & MULT_26(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(69)<=signed(MULT_25(69)(MULT_SIZE-1) & MULT_25(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(69)(MULT_SIZE-1) & MULT_26(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(70)<=signed(MULT_25(70)(MULT_SIZE-1) & MULT_25(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(70)(MULT_SIZE-1) & MULT_26(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(71)<=signed(MULT_25(71)(MULT_SIZE-1) & MULT_25(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(71)(MULT_SIZE-1) & MULT_26(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(72)<=signed(MULT_25(72)(MULT_SIZE-1) & MULT_25(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(72)(MULT_SIZE-1) & MULT_26(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(73)<=signed(MULT_25(73)(MULT_SIZE-1) & MULT_25(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(73)(MULT_SIZE-1) & MULT_26(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(74)<=signed(MULT_25(74)(MULT_SIZE-1) & MULT_25(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(74)(MULT_SIZE-1) & MULT_26(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(75)<=signed(MULT_25(75)(MULT_SIZE-1) & MULT_25(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(75)(MULT_SIZE-1) & MULT_26(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(76)<=signed(MULT_25(76)(MULT_SIZE-1) & MULT_25(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(76)(MULT_SIZE-1) & MULT_26(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(77)<=signed(MULT_25(77)(MULT_SIZE-1) & MULT_25(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(77)(MULT_SIZE-1) & MULT_26(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(78)<=signed(MULT_25(78)(MULT_SIZE-1) & MULT_25(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(78)(MULT_SIZE-1) & MULT_26(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(79)<=signed(MULT_25(79)(MULT_SIZE-1) & MULT_25(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(79)(MULT_SIZE-1) & MULT_26(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(80)<=signed(MULT_25(80)(MULT_SIZE-1) & MULT_25(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(80)(MULT_SIZE-1) & MULT_26(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(81)<=signed(MULT_25(81)(MULT_SIZE-1) & MULT_25(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(81)(MULT_SIZE-1) & MULT_26(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(82)<=signed(MULT_25(82)(MULT_SIZE-1) & MULT_25(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(82)(MULT_SIZE-1) & MULT_26(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13(83)<=signed(MULT_25(83)(MULT_SIZE-1) & MULT_25(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_26(83)(MULT_SIZE-1) & MULT_26(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_14(0)<=signed(MULT_27(0)(MULT_SIZE-1) & MULT_27(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(0)(MULT_SIZE-1) & MULT_28(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(1)<=signed(MULT_27(1)(MULT_SIZE-1) & MULT_27(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(1)(MULT_SIZE-1) & MULT_28(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(2)<=signed(MULT_27(2)(MULT_SIZE-1) & MULT_27(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(2)(MULT_SIZE-1) & MULT_28(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(3)<=signed(MULT_27(3)(MULT_SIZE-1) & MULT_27(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(3)(MULT_SIZE-1) & MULT_28(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(4)<=signed(MULT_27(4)(MULT_SIZE-1) & MULT_27(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(4)(MULT_SIZE-1) & MULT_28(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(5)<=signed(MULT_27(5)(MULT_SIZE-1) & MULT_27(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(5)(MULT_SIZE-1) & MULT_28(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(6)<=signed(MULT_27(6)(MULT_SIZE-1) & MULT_27(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(6)(MULT_SIZE-1) & MULT_28(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(7)<=signed(MULT_27(7)(MULT_SIZE-1) & MULT_27(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(7)(MULT_SIZE-1) & MULT_28(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(8)<=signed(MULT_27(8)(MULT_SIZE-1) & MULT_27(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(8)(MULT_SIZE-1) & MULT_28(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(9)<=signed(MULT_27(9)(MULT_SIZE-1) & MULT_27(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(9)(MULT_SIZE-1) & MULT_28(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(10)<=signed(MULT_27(10)(MULT_SIZE-1) & MULT_27(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(10)(MULT_SIZE-1) & MULT_28(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(11)<=signed(MULT_27(11)(MULT_SIZE-1) & MULT_27(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(11)(MULT_SIZE-1) & MULT_28(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(12)<=signed(MULT_27(12)(MULT_SIZE-1) & MULT_27(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(12)(MULT_SIZE-1) & MULT_28(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(13)<=signed(MULT_27(13)(MULT_SIZE-1) & MULT_27(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(13)(MULT_SIZE-1) & MULT_28(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(14)<=signed(MULT_27(14)(MULT_SIZE-1) & MULT_27(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(14)(MULT_SIZE-1) & MULT_28(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(15)<=signed(MULT_27(15)(MULT_SIZE-1) & MULT_27(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(15)(MULT_SIZE-1) & MULT_28(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(16)<=signed(MULT_27(16)(MULT_SIZE-1) & MULT_27(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(16)(MULT_SIZE-1) & MULT_28(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(17)<=signed(MULT_27(17)(MULT_SIZE-1) & MULT_27(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(17)(MULT_SIZE-1) & MULT_28(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(18)<=signed(MULT_27(18)(MULT_SIZE-1) & MULT_27(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(18)(MULT_SIZE-1) & MULT_28(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(19)<=signed(MULT_27(19)(MULT_SIZE-1) & MULT_27(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(19)(MULT_SIZE-1) & MULT_28(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(20)<=signed(MULT_27(20)(MULT_SIZE-1) & MULT_27(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(20)(MULT_SIZE-1) & MULT_28(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(21)<=signed(MULT_27(21)(MULT_SIZE-1) & MULT_27(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(21)(MULT_SIZE-1) & MULT_28(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(22)<=signed(MULT_27(22)(MULT_SIZE-1) & MULT_27(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(22)(MULT_SIZE-1) & MULT_28(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(23)<=signed(MULT_27(23)(MULT_SIZE-1) & MULT_27(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(23)(MULT_SIZE-1) & MULT_28(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(24)<=signed(MULT_27(24)(MULT_SIZE-1) & MULT_27(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(24)(MULT_SIZE-1) & MULT_28(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(25)<=signed(MULT_27(25)(MULT_SIZE-1) & MULT_27(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(25)(MULT_SIZE-1) & MULT_28(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(26)<=signed(MULT_27(26)(MULT_SIZE-1) & MULT_27(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(26)(MULT_SIZE-1) & MULT_28(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(27)<=signed(MULT_27(27)(MULT_SIZE-1) & MULT_27(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(27)(MULT_SIZE-1) & MULT_28(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(28)<=signed(MULT_27(28)(MULT_SIZE-1) & MULT_27(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(28)(MULT_SIZE-1) & MULT_28(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(29)<=signed(MULT_27(29)(MULT_SIZE-1) & MULT_27(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(29)(MULT_SIZE-1) & MULT_28(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(30)<=signed(MULT_27(30)(MULT_SIZE-1) & MULT_27(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(30)(MULT_SIZE-1) & MULT_28(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(31)<=signed(MULT_27(31)(MULT_SIZE-1) & MULT_27(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(31)(MULT_SIZE-1) & MULT_28(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(32)<=signed(MULT_27(32)(MULT_SIZE-1) & MULT_27(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(32)(MULT_SIZE-1) & MULT_28(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(33)<=signed(MULT_27(33)(MULT_SIZE-1) & MULT_27(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(33)(MULT_SIZE-1) & MULT_28(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(34)<=signed(MULT_27(34)(MULT_SIZE-1) & MULT_27(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(34)(MULT_SIZE-1) & MULT_28(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(35)<=signed(MULT_27(35)(MULT_SIZE-1) & MULT_27(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(35)(MULT_SIZE-1) & MULT_28(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(36)<=signed(MULT_27(36)(MULT_SIZE-1) & MULT_27(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(36)(MULT_SIZE-1) & MULT_28(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(37)<=signed(MULT_27(37)(MULT_SIZE-1) & MULT_27(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(37)(MULT_SIZE-1) & MULT_28(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(38)<=signed(MULT_27(38)(MULT_SIZE-1) & MULT_27(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(38)(MULT_SIZE-1) & MULT_28(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(39)<=signed(MULT_27(39)(MULT_SIZE-1) & MULT_27(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(39)(MULT_SIZE-1) & MULT_28(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(40)<=signed(MULT_27(40)(MULT_SIZE-1) & MULT_27(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(40)(MULT_SIZE-1) & MULT_28(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(41)<=signed(MULT_27(41)(MULT_SIZE-1) & MULT_27(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(41)(MULT_SIZE-1) & MULT_28(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(42)<=signed(MULT_27(42)(MULT_SIZE-1) & MULT_27(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(42)(MULT_SIZE-1) & MULT_28(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(43)<=signed(MULT_27(43)(MULT_SIZE-1) & MULT_27(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(43)(MULT_SIZE-1) & MULT_28(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(44)<=signed(MULT_27(44)(MULT_SIZE-1) & MULT_27(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(44)(MULT_SIZE-1) & MULT_28(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(45)<=signed(MULT_27(45)(MULT_SIZE-1) & MULT_27(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(45)(MULT_SIZE-1) & MULT_28(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(46)<=signed(MULT_27(46)(MULT_SIZE-1) & MULT_27(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(46)(MULT_SIZE-1) & MULT_28(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(47)<=signed(MULT_27(47)(MULT_SIZE-1) & MULT_27(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(47)(MULT_SIZE-1) & MULT_28(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(48)<=signed(MULT_27(48)(MULT_SIZE-1) & MULT_27(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(48)(MULT_SIZE-1) & MULT_28(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(49)<=signed(MULT_27(49)(MULT_SIZE-1) & MULT_27(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(49)(MULT_SIZE-1) & MULT_28(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(50)<=signed(MULT_27(50)(MULT_SIZE-1) & MULT_27(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(50)(MULT_SIZE-1) & MULT_28(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(51)<=signed(MULT_27(51)(MULT_SIZE-1) & MULT_27(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(51)(MULT_SIZE-1) & MULT_28(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(52)<=signed(MULT_27(52)(MULT_SIZE-1) & MULT_27(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(52)(MULT_SIZE-1) & MULT_28(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(53)<=signed(MULT_27(53)(MULT_SIZE-1) & MULT_27(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(53)(MULT_SIZE-1) & MULT_28(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(54)<=signed(MULT_27(54)(MULT_SIZE-1) & MULT_27(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(54)(MULT_SIZE-1) & MULT_28(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(55)<=signed(MULT_27(55)(MULT_SIZE-1) & MULT_27(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(55)(MULT_SIZE-1) & MULT_28(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(56)<=signed(MULT_27(56)(MULT_SIZE-1) & MULT_27(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(56)(MULT_SIZE-1) & MULT_28(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(57)<=signed(MULT_27(57)(MULT_SIZE-1) & MULT_27(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(57)(MULT_SIZE-1) & MULT_28(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(58)<=signed(MULT_27(58)(MULT_SIZE-1) & MULT_27(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(58)(MULT_SIZE-1) & MULT_28(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(59)<=signed(MULT_27(59)(MULT_SIZE-1) & MULT_27(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(59)(MULT_SIZE-1) & MULT_28(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(60)<=signed(MULT_27(60)(MULT_SIZE-1) & MULT_27(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(60)(MULT_SIZE-1) & MULT_28(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(61)<=signed(MULT_27(61)(MULT_SIZE-1) & MULT_27(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(61)(MULT_SIZE-1) & MULT_28(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(62)<=signed(MULT_27(62)(MULT_SIZE-1) & MULT_27(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(62)(MULT_SIZE-1) & MULT_28(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(63)<=signed(MULT_27(63)(MULT_SIZE-1) & MULT_27(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(63)(MULT_SIZE-1) & MULT_28(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(64)<=signed(MULT_27(64)(MULT_SIZE-1) & MULT_27(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(64)(MULT_SIZE-1) & MULT_28(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(65)<=signed(MULT_27(65)(MULT_SIZE-1) & MULT_27(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(65)(MULT_SIZE-1) & MULT_28(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(66)<=signed(MULT_27(66)(MULT_SIZE-1) & MULT_27(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(66)(MULT_SIZE-1) & MULT_28(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(67)<=signed(MULT_27(67)(MULT_SIZE-1) & MULT_27(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(67)(MULT_SIZE-1) & MULT_28(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(68)<=signed(MULT_27(68)(MULT_SIZE-1) & MULT_27(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(68)(MULT_SIZE-1) & MULT_28(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(69)<=signed(MULT_27(69)(MULT_SIZE-1) & MULT_27(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(69)(MULT_SIZE-1) & MULT_28(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(70)<=signed(MULT_27(70)(MULT_SIZE-1) & MULT_27(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(70)(MULT_SIZE-1) & MULT_28(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(71)<=signed(MULT_27(71)(MULT_SIZE-1) & MULT_27(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(71)(MULT_SIZE-1) & MULT_28(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(72)<=signed(MULT_27(72)(MULT_SIZE-1) & MULT_27(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(72)(MULT_SIZE-1) & MULT_28(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(73)<=signed(MULT_27(73)(MULT_SIZE-1) & MULT_27(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(73)(MULT_SIZE-1) & MULT_28(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(74)<=signed(MULT_27(74)(MULT_SIZE-1) & MULT_27(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(74)(MULT_SIZE-1) & MULT_28(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(75)<=signed(MULT_27(75)(MULT_SIZE-1) & MULT_27(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(75)(MULT_SIZE-1) & MULT_28(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(76)<=signed(MULT_27(76)(MULT_SIZE-1) & MULT_27(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(76)(MULT_SIZE-1) & MULT_28(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(77)<=signed(MULT_27(77)(MULT_SIZE-1) & MULT_27(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(77)(MULT_SIZE-1) & MULT_28(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(78)<=signed(MULT_27(78)(MULT_SIZE-1) & MULT_27(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(78)(MULT_SIZE-1) & MULT_28(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(79)<=signed(MULT_27(79)(MULT_SIZE-1) & MULT_27(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(79)(MULT_SIZE-1) & MULT_28(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(80)<=signed(MULT_27(80)(MULT_SIZE-1) & MULT_27(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(80)(MULT_SIZE-1) & MULT_28(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(81)<=signed(MULT_27(81)(MULT_SIZE-1) & MULT_27(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(81)(MULT_SIZE-1) & MULT_28(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(82)<=signed(MULT_27(82)(MULT_SIZE-1) & MULT_27(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(82)(MULT_SIZE-1) & MULT_28(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14(83)<=signed(MULT_27(83)(MULT_SIZE-1) & MULT_27(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_28(83)(MULT_SIZE-1) & MULT_28(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_15(0)<=signed(MULT_29(0)(MULT_SIZE-1) & MULT_29(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(0)(MULT_SIZE-1) & MULT_30(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(1)<=signed(MULT_29(1)(MULT_SIZE-1) & MULT_29(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(1)(MULT_SIZE-1) & MULT_30(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(2)<=signed(MULT_29(2)(MULT_SIZE-1) & MULT_29(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(2)(MULT_SIZE-1) & MULT_30(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(3)<=signed(MULT_29(3)(MULT_SIZE-1) & MULT_29(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(3)(MULT_SIZE-1) & MULT_30(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(4)<=signed(MULT_29(4)(MULT_SIZE-1) & MULT_29(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(4)(MULT_SIZE-1) & MULT_30(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(5)<=signed(MULT_29(5)(MULT_SIZE-1) & MULT_29(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(5)(MULT_SIZE-1) & MULT_30(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(6)<=signed(MULT_29(6)(MULT_SIZE-1) & MULT_29(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(6)(MULT_SIZE-1) & MULT_30(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(7)<=signed(MULT_29(7)(MULT_SIZE-1) & MULT_29(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(7)(MULT_SIZE-1) & MULT_30(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(8)<=signed(MULT_29(8)(MULT_SIZE-1) & MULT_29(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(8)(MULT_SIZE-1) & MULT_30(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(9)<=signed(MULT_29(9)(MULT_SIZE-1) & MULT_29(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(9)(MULT_SIZE-1) & MULT_30(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(10)<=signed(MULT_29(10)(MULT_SIZE-1) & MULT_29(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(10)(MULT_SIZE-1) & MULT_30(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(11)<=signed(MULT_29(11)(MULT_SIZE-1) & MULT_29(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(11)(MULT_SIZE-1) & MULT_30(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(12)<=signed(MULT_29(12)(MULT_SIZE-1) & MULT_29(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(12)(MULT_SIZE-1) & MULT_30(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(13)<=signed(MULT_29(13)(MULT_SIZE-1) & MULT_29(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(13)(MULT_SIZE-1) & MULT_30(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(14)<=signed(MULT_29(14)(MULT_SIZE-1) & MULT_29(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(14)(MULT_SIZE-1) & MULT_30(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(15)<=signed(MULT_29(15)(MULT_SIZE-1) & MULT_29(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(15)(MULT_SIZE-1) & MULT_30(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(16)<=signed(MULT_29(16)(MULT_SIZE-1) & MULT_29(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(16)(MULT_SIZE-1) & MULT_30(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(17)<=signed(MULT_29(17)(MULT_SIZE-1) & MULT_29(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(17)(MULT_SIZE-1) & MULT_30(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(18)<=signed(MULT_29(18)(MULT_SIZE-1) & MULT_29(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(18)(MULT_SIZE-1) & MULT_30(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(19)<=signed(MULT_29(19)(MULT_SIZE-1) & MULT_29(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(19)(MULT_SIZE-1) & MULT_30(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(20)<=signed(MULT_29(20)(MULT_SIZE-1) & MULT_29(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(20)(MULT_SIZE-1) & MULT_30(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(21)<=signed(MULT_29(21)(MULT_SIZE-1) & MULT_29(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(21)(MULT_SIZE-1) & MULT_30(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(22)<=signed(MULT_29(22)(MULT_SIZE-1) & MULT_29(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(22)(MULT_SIZE-1) & MULT_30(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(23)<=signed(MULT_29(23)(MULT_SIZE-1) & MULT_29(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(23)(MULT_SIZE-1) & MULT_30(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(24)<=signed(MULT_29(24)(MULT_SIZE-1) & MULT_29(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(24)(MULT_SIZE-1) & MULT_30(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(25)<=signed(MULT_29(25)(MULT_SIZE-1) & MULT_29(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(25)(MULT_SIZE-1) & MULT_30(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(26)<=signed(MULT_29(26)(MULT_SIZE-1) & MULT_29(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(26)(MULT_SIZE-1) & MULT_30(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(27)<=signed(MULT_29(27)(MULT_SIZE-1) & MULT_29(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(27)(MULT_SIZE-1) & MULT_30(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(28)<=signed(MULT_29(28)(MULT_SIZE-1) & MULT_29(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(28)(MULT_SIZE-1) & MULT_30(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(29)<=signed(MULT_29(29)(MULT_SIZE-1) & MULT_29(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(29)(MULT_SIZE-1) & MULT_30(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(30)<=signed(MULT_29(30)(MULT_SIZE-1) & MULT_29(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(30)(MULT_SIZE-1) & MULT_30(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(31)<=signed(MULT_29(31)(MULT_SIZE-1) & MULT_29(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(31)(MULT_SIZE-1) & MULT_30(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(32)<=signed(MULT_29(32)(MULT_SIZE-1) & MULT_29(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(32)(MULT_SIZE-1) & MULT_30(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(33)<=signed(MULT_29(33)(MULT_SIZE-1) & MULT_29(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(33)(MULT_SIZE-1) & MULT_30(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(34)<=signed(MULT_29(34)(MULT_SIZE-1) & MULT_29(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(34)(MULT_SIZE-1) & MULT_30(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(35)<=signed(MULT_29(35)(MULT_SIZE-1) & MULT_29(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(35)(MULT_SIZE-1) & MULT_30(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(36)<=signed(MULT_29(36)(MULT_SIZE-1) & MULT_29(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(36)(MULT_SIZE-1) & MULT_30(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(37)<=signed(MULT_29(37)(MULT_SIZE-1) & MULT_29(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(37)(MULT_SIZE-1) & MULT_30(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(38)<=signed(MULT_29(38)(MULT_SIZE-1) & MULT_29(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(38)(MULT_SIZE-1) & MULT_30(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(39)<=signed(MULT_29(39)(MULT_SIZE-1) & MULT_29(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(39)(MULT_SIZE-1) & MULT_30(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(40)<=signed(MULT_29(40)(MULT_SIZE-1) & MULT_29(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(40)(MULT_SIZE-1) & MULT_30(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(41)<=signed(MULT_29(41)(MULT_SIZE-1) & MULT_29(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(41)(MULT_SIZE-1) & MULT_30(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(42)<=signed(MULT_29(42)(MULT_SIZE-1) & MULT_29(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(42)(MULT_SIZE-1) & MULT_30(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(43)<=signed(MULT_29(43)(MULT_SIZE-1) & MULT_29(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(43)(MULT_SIZE-1) & MULT_30(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(44)<=signed(MULT_29(44)(MULT_SIZE-1) & MULT_29(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(44)(MULT_SIZE-1) & MULT_30(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(45)<=signed(MULT_29(45)(MULT_SIZE-1) & MULT_29(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(45)(MULT_SIZE-1) & MULT_30(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(46)<=signed(MULT_29(46)(MULT_SIZE-1) & MULT_29(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(46)(MULT_SIZE-1) & MULT_30(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(47)<=signed(MULT_29(47)(MULT_SIZE-1) & MULT_29(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(47)(MULT_SIZE-1) & MULT_30(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(48)<=signed(MULT_29(48)(MULT_SIZE-1) & MULT_29(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(48)(MULT_SIZE-1) & MULT_30(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(49)<=signed(MULT_29(49)(MULT_SIZE-1) & MULT_29(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(49)(MULT_SIZE-1) & MULT_30(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(50)<=signed(MULT_29(50)(MULT_SIZE-1) & MULT_29(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(50)(MULT_SIZE-1) & MULT_30(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(51)<=signed(MULT_29(51)(MULT_SIZE-1) & MULT_29(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(51)(MULT_SIZE-1) & MULT_30(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(52)<=signed(MULT_29(52)(MULT_SIZE-1) & MULT_29(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(52)(MULT_SIZE-1) & MULT_30(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(53)<=signed(MULT_29(53)(MULT_SIZE-1) & MULT_29(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(53)(MULT_SIZE-1) & MULT_30(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(54)<=signed(MULT_29(54)(MULT_SIZE-1) & MULT_29(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(54)(MULT_SIZE-1) & MULT_30(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(55)<=signed(MULT_29(55)(MULT_SIZE-1) & MULT_29(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(55)(MULT_SIZE-1) & MULT_30(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(56)<=signed(MULT_29(56)(MULT_SIZE-1) & MULT_29(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(56)(MULT_SIZE-1) & MULT_30(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(57)<=signed(MULT_29(57)(MULT_SIZE-1) & MULT_29(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(57)(MULT_SIZE-1) & MULT_30(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(58)<=signed(MULT_29(58)(MULT_SIZE-1) & MULT_29(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(58)(MULT_SIZE-1) & MULT_30(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(59)<=signed(MULT_29(59)(MULT_SIZE-1) & MULT_29(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(59)(MULT_SIZE-1) & MULT_30(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(60)<=signed(MULT_29(60)(MULT_SIZE-1) & MULT_29(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(60)(MULT_SIZE-1) & MULT_30(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(61)<=signed(MULT_29(61)(MULT_SIZE-1) & MULT_29(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(61)(MULT_SIZE-1) & MULT_30(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(62)<=signed(MULT_29(62)(MULT_SIZE-1) & MULT_29(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(62)(MULT_SIZE-1) & MULT_30(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(63)<=signed(MULT_29(63)(MULT_SIZE-1) & MULT_29(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(63)(MULT_SIZE-1) & MULT_30(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(64)<=signed(MULT_29(64)(MULT_SIZE-1) & MULT_29(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(64)(MULT_SIZE-1) & MULT_30(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(65)<=signed(MULT_29(65)(MULT_SIZE-1) & MULT_29(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(65)(MULT_SIZE-1) & MULT_30(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(66)<=signed(MULT_29(66)(MULT_SIZE-1) & MULT_29(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(66)(MULT_SIZE-1) & MULT_30(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(67)<=signed(MULT_29(67)(MULT_SIZE-1) & MULT_29(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(67)(MULT_SIZE-1) & MULT_30(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(68)<=signed(MULT_29(68)(MULT_SIZE-1) & MULT_29(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(68)(MULT_SIZE-1) & MULT_30(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(69)<=signed(MULT_29(69)(MULT_SIZE-1) & MULT_29(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(69)(MULT_SIZE-1) & MULT_30(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(70)<=signed(MULT_29(70)(MULT_SIZE-1) & MULT_29(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(70)(MULT_SIZE-1) & MULT_30(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(71)<=signed(MULT_29(71)(MULT_SIZE-1) & MULT_29(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(71)(MULT_SIZE-1) & MULT_30(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(72)<=signed(MULT_29(72)(MULT_SIZE-1) & MULT_29(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(72)(MULT_SIZE-1) & MULT_30(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(73)<=signed(MULT_29(73)(MULT_SIZE-1) & MULT_29(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(73)(MULT_SIZE-1) & MULT_30(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(74)<=signed(MULT_29(74)(MULT_SIZE-1) & MULT_29(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(74)(MULT_SIZE-1) & MULT_30(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(75)<=signed(MULT_29(75)(MULT_SIZE-1) & MULT_29(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(75)(MULT_SIZE-1) & MULT_30(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(76)<=signed(MULT_29(76)(MULT_SIZE-1) & MULT_29(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(76)(MULT_SIZE-1) & MULT_30(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(77)<=signed(MULT_29(77)(MULT_SIZE-1) & MULT_29(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(77)(MULT_SIZE-1) & MULT_30(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(78)<=signed(MULT_29(78)(MULT_SIZE-1) & MULT_29(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(78)(MULT_SIZE-1) & MULT_30(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(79)<=signed(MULT_29(79)(MULT_SIZE-1) & MULT_29(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(79)(MULT_SIZE-1) & MULT_30(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(80)<=signed(MULT_29(80)(MULT_SIZE-1) & MULT_29(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(80)(MULT_SIZE-1) & MULT_30(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(81)<=signed(MULT_29(81)(MULT_SIZE-1) & MULT_29(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(81)(MULT_SIZE-1) & MULT_30(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(82)<=signed(MULT_29(82)(MULT_SIZE-1) & MULT_29(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(82)(MULT_SIZE-1) & MULT_30(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15(83)<=signed(MULT_29(83)(MULT_SIZE-1) & MULT_29(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_30(83)(MULT_SIZE-1) & MULT_30(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_16(0)<=signed(MULT_31(0)(MULT_SIZE-1) & MULT_31(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(0)(MULT_SIZE-1) & MULT_32(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(1)<=signed(MULT_31(1)(MULT_SIZE-1) & MULT_31(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(1)(MULT_SIZE-1) & MULT_32(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(2)<=signed(MULT_31(2)(MULT_SIZE-1) & MULT_31(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(2)(MULT_SIZE-1) & MULT_32(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(3)<=signed(MULT_31(3)(MULT_SIZE-1) & MULT_31(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(3)(MULT_SIZE-1) & MULT_32(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(4)<=signed(MULT_31(4)(MULT_SIZE-1) & MULT_31(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(4)(MULT_SIZE-1) & MULT_32(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(5)<=signed(MULT_31(5)(MULT_SIZE-1) & MULT_31(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(5)(MULT_SIZE-1) & MULT_32(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(6)<=signed(MULT_31(6)(MULT_SIZE-1) & MULT_31(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(6)(MULT_SIZE-1) & MULT_32(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(7)<=signed(MULT_31(7)(MULT_SIZE-1) & MULT_31(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(7)(MULT_SIZE-1) & MULT_32(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(8)<=signed(MULT_31(8)(MULT_SIZE-1) & MULT_31(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(8)(MULT_SIZE-1) & MULT_32(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(9)<=signed(MULT_31(9)(MULT_SIZE-1) & MULT_31(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(9)(MULT_SIZE-1) & MULT_32(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(10)<=signed(MULT_31(10)(MULT_SIZE-1) & MULT_31(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(10)(MULT_SIZE-1) & MULT_32(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(11)<=signed(MULT_31(11)(MULT_SIZE-1) & MULT_31(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(11)(MULT_SIZE-1) & MULT_32(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(12)<=signed(MULT_31(12)(MULT_SIZE-1) & MULT_31(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(12)(MULT_SIZE-1) & MULT_32(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(13)<=signed(MULT_31(13)(MULT_SIZE-1) & MULT_31(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(13)(MULT_SIZE-1) & MULT_32(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(14)<=signed(MULT_31(14)(MULT_SIZE-1) & MULT_31(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(14)(MULT_SIZE-1) & MULT_32(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(15)<=signed(MULT_31(15)(MULT_SIZE-1) & MULT_31(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(15)(MULT_SIZE-1) & MULT_32(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(16)<=signed(MULT_31(16)(MULT_SIZE-1) & MULT_31(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(16)(MULT_SIZE-1) & MULT_32(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(17)<=signed(MULT_31(17)(MULT_SIZE-1) & MULT_31(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(17)(MULT_SIZE-1) & MULT_32(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(18)<=signed(MULT_31(18)(MULT_SIZE-1) & MULT_31(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(18)(MULT_SIZE-1) & MULT_32(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(19)<=signed(MULT_31(19)(MULT_SIZE-1) & MULT_31(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(19)(MULT_SIZE-1) & MULT_32(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(20)<=signed(MULT_31(20)(MULT_SIZE-1) & MULT_31(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(20)(MULT_SIZE-1) & MULT_32(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(21)<=signed(MULT_31(21)(MULT_SIZE-1) & MULT_31(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(21)(MULT_SIZE-1) & MULT_32(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(22)<=signed(MULT_31(22)(MULT_SIZE-1) & MULT_31(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(22)(MULT_SIZE-1) & MULT_32(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(23)<=signed(MULT_31(23)(MULT_SIZE-1) & MULT_31(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(23)(MULT_SIZE-1) & MULT_32(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(24)<=signed(MULT_31(24)(MULT_SIZE-1) & MULT_31(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(24)(MULT_SIZE-1) & MULT_32(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(25)<=signed(MULT_31(25)(MULT_SIZE-1) & MULT_31(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(25)(MULT_SIZE-1) & MULT_32(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(26)<=signed(MULT_31(26)(MULT_SIZE-1) & MULT_31(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(26)(MULT_SIZE-1) & MULT_32(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(27)<=signed(MULT_31(27)(MULT_SIZE-1) & MULT_31(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(27)(MULT_SIZE-1) & MULT_32(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(28)<=signed(MULT_31(28)(MULT_SIZE-1) & MULT_31(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(28)(MULT_SIZE-1) & MULT_32(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(29)<=signed(MULT_31(29)(MULT_SIZE-1) & MULT_31(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(29)(MULT_SIZE-1) & MULT_32(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(30)<=signed(MULT_31(30)(MULT_SIZE-1) & MULT_31(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(30)(MULT_SIZE-1) & MULT_32(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(31)<=signed(MULT_31(31)(MULT_SIZE-1) & MULT_31(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(31)(MULT_SIZE-1) & MULT_32(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(32)<=signed(MULT_31(32)(MULT_SIZE-1) & MULT_31(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(32)(MULT_SIZE-1) & MULT_32(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(33)<=signed(MULT_31(33)(MULT_SIZE-1) & MULT_31(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(33)(MULT_SIZE-1) & MULT_32(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(34)<=signed(MULT_31(34)(MULT_SIZE-1) & MULT_31(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(34)(MULT_SIZE-1) & MULT_32(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(35)<=signed(MULT_31(35)(MULT_SIZE-1) & MULT_31(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(35)(MULT_SIZE-1) & MULT_32(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(36)<=signed(MULT_31(36)(MULT_SIZE-1) & MULT_31(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(36)(MULT_SIZE-1) & MULT_32(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(37)<=signed(MULT_31(37)(MULT_SIZE-1) & MULT_31(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(37)(MULT_SIZE-1) & MULT_32(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(38)<=signed(MULT_31(38)(MULT_SIZE-1) & MULT_31(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(38)(MULT_SIZE-1) & MULT_32(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(39)<=signed(MULT_31(39)(MULT_SIZE-1) & MULT_31(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(39)(MULT_SIZE-1) & MULT_32(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(40)<=signed(MULT_31(40)(MULT_SIZE-1) & MULT_31(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(40)(MULT_SIZE-1) & MULT_32(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(41)<=signed(MULT_31(41)(MULT_SIZE-1) & MULT_31(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(41)(MULT_SIZE-1) & MULT_32(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(42)<=signed(MULT_31(42)(MULT_SIZE-1) & MULT_31(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(42)(MULT_SIZE-1) & MULT_32(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(43)<=signed(MULT_31(43)(MULT_SIZE-1) & MULT_31(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(43)(MULT_SIZE-1) & MULT_32(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(44)<=signed(MULT_31(44)(MULT_SIZE-1) & MULT_31(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(44)(MULT_SIZE-1) & MULT_32(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(45)<=signed(MULT_31(45)(MULT_SIZE-1) & MULT_31(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(45)(MULT_SIZE-1) & MULT_32(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(46)<=signed(MULT_31(46)(MULT_SIZE-1) & MULT_31(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(46)(MULT_SIZE-1) & MULT_32(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(47)<=signed(MULT_31(47)(MULT_SIZE-1) & MULT_31(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(47)(MULT_SIZE-1) & MULT_32(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(48)<=signed(MULT_31(48)(MULT_SIZE-1) & MULT_31(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(48)(MULT_SIZE-1) & MULT_32(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(49)<=signed(MULT_31(49)(MULT_SIZE-1) & MULT_31(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(49)(MULT_SIZE-1) & MULT_32(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(50)<=signed(MULT_31(50)(MULT_SIZE-1) & MULT_31(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(50)(MULT_SIZE-1) & MULT_32(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(51)<=signed(MULT_31(51)(MULT_SIZE-1) & MULT_31(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(51)(MULT_SIZE-1) & MULT_32(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(52)<=signed(MULT_31(52)(MULT_SIZE-1) & MULT_31(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(52)(MULT_SIZE-1) & MULT_32(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(53)<=signed(MULT_31(53)(MULT_SIZE-1) & MULT_31(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(53)(MULT_SIZE-1) & MULT_32(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(54)<=signed(MULT_31(54)(MULT_SIZE-1) & MULT_31(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(54)(MULT_SIZE-1) & MULT_32(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(55)<=signed(MULT_31(55)(MULT_SIZE-1) & MULT_31(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(55)(MULT_SIZE-1) & MULT_32(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(56)<=signed(MULT_31(56)(MULT_SIZE-1) & MULT_31(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(56)(MULT_SIZE-1) & MULT_32(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(57)<=signed(MULT_31(57)(MULT_SIZE-1) & MULT_31(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(57)(MULT_SIZE-1) & MULT_32(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(58)<=signed(MULT_31(58)(MULT_SIZE-1) & MULT_31(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(58)(MULT_SIZE-1) & MULT_32(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(59)<=signed(MULT_31(59)(MULT_SIZE-1) & MULT_31(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(59)(MULT_SIZE-1) & MULT_32(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(60)<=signed(MULT_31(60)(MULT_SIZE-1) & MULT_31(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(60)(MULT_SIZE-1) & MULT_32(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(61)<=signed(MULT_31(61)(MULT_SIZE-1) & MULT_31(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(61)(MULT_SIZE-1) & MULT_32(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(62)<=signed(MULT_31(62)(MULT_SIZE-1) & MULT_31(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(62)(MULT_SIZE-1) & MULT_32(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(63)<=signed(MULT_31(63)(MULT_SIZE-1) & MULT_31(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(63)(MULT_SIZE-1) & MULT_32(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(64)<=signed(MULT_31(64)(MULT_SIZE-1) & MULT_31(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(64)(MULT_SIZE-1) & MULT_32(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(65)<=signed(MULT_31(65)(MULT_SIZE-1) & MULT_31(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(65)(MULT_SIZE-1) & MULT_32(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(66)<=signed(MULT_31(66)(MULT_SIZE-1) & MULT_31(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(66)(MULT_SIZE-1) & MULT_32(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(67)<=signed(MULT_31(67)(MULT_SIZE-1) & MULT_31(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(67)(MULT_SIZE-1) & MULT_32(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(68)<=signed(MULT_31(68)(MULT_SIZE-1) & MULT_31(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(68)(MULT_SIZE-1) & MULT_32(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(69)<=signed(MULT_31(69)(MULT_SIZE-1) & MULT_31(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(69)(MULT_SIZE-1) & MULT_32(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(70)<=signed(MULT_31(70)(MULT_SIZE-1) & MULT_31(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(70)(MULT_SIZE-1) & MULT_32(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(71)<=signed(MULT_31(71)(MULT_SIZE-1) & MULT_31(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(71)(MULT_SIZE-1) & MULT_32(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(72)<=signed(MULT_31(72)(MULT_SIZE-1) & MULT_31(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(72)(MULT_SIZE-1) & MULT_32(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(73)<=signed(MULT_31(73)(MULT_SIZE-1) & MULT_31(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(73)(MULT_SIZE-1) & MULT_32(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(74)<=signed(MULT_31(74)(MULT_SIZE-1) & MULT_31(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(74)(MULT_SIZE-1) & MULT_32(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(75)<=signed(MULT_31(75)(MULT_SIZE-1) & MULT_31(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(75)(MULT_SIZE-1) & MULT_32(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(76)<=signed(MULT_31(76)(MULT_SIZE-1) & MULT_31(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(76)(MULT_SIZE-1) & MULT_32(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(77)<=signed(MULT_31(77)(MULT_SIZE-1) & MULT_31(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(77)(MULT_SIZE-1) & MULT_32(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(78)<=signed(MULT_31(78)(MULT_SIZE-1) & MULT_31(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(78)(MULT_SIZE-1) & MULT_32(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(79)<=signed(MULT_31(79)(MULT_SIZE-1) & MULT_31(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(79)(MULT_SIZE-1) & MULT_32(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(80)<=signed(MULT_31(80)(MULT_SIZE-1) & MULT_31(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(80)(MULT_SIZE-1) & MULT_32(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(81)<=signed(MULT_31(81)(MULT_SIZE-1) & MULT_31(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(81)(MULT_SIZE-1) & MULT_32(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(82)<=signed(MULT_31(82)(MULT_SIZE-1) & MULT_31(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(82)(MULT_SIZE-1) & MULT_32(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16(83)<=signed(MULT_31(83)(MULT_SIZE-1) & MULT_31(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_32(83)(MULT_SIZE-1) & MULT_32(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_17(0)<=signed(MULT_33(0)(MULT_SIZE-1) & MULT_33(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(0)(MULT_SIZE-1) & MULT_34(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(1)<=signed(MULT_33(1)(MULT_SIZE-1) & MULT_33(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(1)(MULT_SIZE-1) & MULT_34(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(2)<=signed(MULT_33(2)(MULT_SIZE-1) & MULT_33(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(2)(MULT_SIZE-1) & MULT_34(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(3)<=signed(MULT_33(3)(MULT_SIZE-1) & MULT_33(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(3)(MULT_SIZE-1) & MULT_34(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(4)<=signed(MULT_33(4)(MULT_SIZE-1) & MULT_33(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(4)(MULT_SIZE-1) & MULT_34(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(5)<=signed(MULT_33(5)(MULT_SIZE-1) & MULT_33(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(5)(MULT_SIZE-1) & MULT_34(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(6)<=signed(MULT_33(6)(MULT_SIZE-1) & MULT_33(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(6)(MULT_SIZE-1) & MULT_34(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(7)<=signed(MULT_33(7)(MULT_SIZE-1) & MULT_33(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(7)(MULT_SIZE-1) & MULT_34(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(8)<=signed(MULT_33(8)(MULT_SIZE-1) & MULT_33(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(8)(MULT_SIZE-1) & MULT_34(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(9)<=signed(MULT_33(9)(MULT_SIZE-1) & MULT_33(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(9)(MULT_SIZE-1) & MULT_34(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(10)<=signed(MULT_33(10)(MULT_SIZE-1) & MULT_33(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(10)(MULT_SIZE-1) & MULT_34(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(11)<=signed(MULT_33(11)(MULT_SIZE-1) & MULT_33(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(11)(MULT_SIZE-1) & MULT_34(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(12)<=signed(MULT_33(12)(MULT_SIZE-1) & MULT_33(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(12)(MULT_SIZE-1) & MULT_34(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(13)<=signed(MULT_33(13)(MULT_SIZE-1) & MULT_33(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(13)(MULT_SIZE-1) & MULT_34(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(14)<=signed(MULT_33(14)(MULT_SIZE-1) & MULT_33(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(14)(MULT_SIZE-1) & MULT_34(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(15)<=signed(MULT_33(15)(MULT_SIZE-1) & MULT_33(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(15)(MULT_SIZE-1) & MULT_34(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(16)<=signed(MULT_33(16)(MULT_SIZE-1) & MULT_33(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(16)(MULT_SIZE-1) & MULT_34(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(17)<=signed(MULT_33(17)(MULT_SIZE-1) & MULT_33(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(17)(MULT_SIZE-1) & MULT_34(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(18)<=signed(MULT_33(18)(MULT_SIZE-1) & MULT_33(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(18)(MULT_SIZE-1) & MULT_34(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(19)<=signed(MULT_33(19)(MULT_SIZE-1) & MULT_33(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(19)(MULT_SIZE-1) & MULT_34(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(20)<=signed(MULT_33(20)(MULT_SIZE-1) & MULT_33(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(20)(MULT_SIZE-1) & MULT_34(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(21)<=signed(MULT_33(21)(MULT_SIZE-1) & MULT_33(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(21)(MULT_SIZE-1) & MULT_34(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(22)<=signed(MULT_33(22)(MULT_SIZE-1) & MULT_33(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(22)(MULT_SIZE-1) & MULT_34(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(23)<=signed(MULT_33(23)(MULT_SIZE-1) & MULT_33(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(23)(MULT_SIZE-1) & MULT_34(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(24)<=signed(MULT_33(24)(MULT_SIZE-1) & MULT_33(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(24)(MULT_SIZE-1) & MULT_34(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(25)<=signed(MULT_33(25)(MULT_SIZE-1) & MULT_33(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(25)(MULT_SIZE-1) & MULT_34(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(26)<=signed(MULT_33(26)(MULT_SIZE-1) & MULT_33(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(26)(MULT_SIZE-1) & MULT_34(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(27)<=signed(MULT_33(27)(MULT_SIZE-1) & MULT_33(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(27)(MULT_SIZE-1) & MULT_34(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(28)<=signed(MULT_33(28)(MULT_SIZE-1) & MULT_33(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(28)(MULT_SIZE-1) & MULT_34(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(29)<=signed(MULT_33(29)(MULT_SIZE-1) & MULT_33(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(29)(MULT_SIZE-1) & MULT_34(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(30)<=signed(MULT_33(30)(MULT_SIZE-1) & MULT_33(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(30)(MULT_SIZE-1) & MULT_34(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(31)<=signed(MULT_33(31)(MULT_SIZE-1) & MULT_33(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(31)(MULT_SIZE-1) & MULT_34(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(32)<=signed(MULT_33(32)(MULT_SIZE-1) & MULT_33(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(32)(MULT_SIZE-1) & MULT_34(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(33)<=signed(MULT_33(33)(MULT_SIZE-1) & MULT_33(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(33)(MULT_SIZE-1) & MULT_34(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(34)<=signed(MULT_33(34)(MULT_SIZE-1) & MULT_33(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(34)(MULT_SIZE-1) & MULT_34(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(35)<=signed(MULT_33(35)(MULT_SIZE-1) & MULT_33(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(35)(MULT_SIZE-1) & MULT_34(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(36)<=signed(MULT_33(36)(MULT_SIZE-1) & MULT_33(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(36)(MULT_SIZE-1) & MULT_34(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(37)<=signed(MULT_33(37)(MULT_SIZE-1) & MULT_33(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(37)(MULT_SIZE-1) & MULT_34(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(38)<=signed(MULT_33(38)(MULT_SIZE-1) & MULT_33(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(38)(MULT_SIZE-1) & MULT_34(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(39)<=signed(MULT_33(39)(MULT_SIZE-1) & MULT_33(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(39)(MULT_SIZE-1) & MULT_34(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(40)<=signed(MULT_33(40)(MULT_SIZE-1) & MULT_33(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(40)(MULT_SIZE-1) & MULT_34(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(41)<=signed(MULT_33(41)(MULT_SIZE-1) & MULT_33(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(41)(MULT_SIZE-1) & MULT_34(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(42)<=signed(MULT_33(42)(MULT_SIZE-1) & MULT_33(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(42)(MULT_SIZE-1) & MULT_34(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(43)<=signed(MULT_33(43)(MULT_SIZE-1) & MULT_33(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(43)(MULT_SIZE-1) & MULT_34(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(44)<=signed(MULT_33(44)(MULT_SIZE-1) & MULT_33(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(44)(MULT_SIZE-1) & MULT_34(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(45)<=signed(MULT_33(45)(MULT_SIZE-1) & MULT_33(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(45)(MULT_SIZE-1) & MULT_34(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(46)<=signed(MULT_33(46)(MULT_SIZE-1) & MULT_33(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(46)(MULT_SIZE-1) & MULT_34(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(47)<=signed(MULT_33(47)(MULT_SIZE-1) & MULT_33(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(47)(MULT_SIZE-1) & MULT_34(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(48)<=signed(MULT_33(48)(MULT_SIZE-1) & MULT_33(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(48)(MULT_SIZE-1) & MULT_34(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(49)<=signed(MULT_33(49)(MULT_SIZE-1) & MULT_33(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(49)(MULT_SIZE-1) & MULT_34(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(50)<=signed(MULT_33(50)(MULT_SIZE-1) & MULT_33(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(50)(MULT_SIZE-1) & MULT_34(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(51)<=signed(MULT_33(51)(MULT_SIZE-1) & MULT_33(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(51)(MULT_SIZE-1) & MULT_34(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(52)<=signed(MULT_33(52)(MULT_SIZE-1) & MULT_33(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(52)(MULT_SIZE-1) & MULT_34(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(53)<=signed(MULT_33(53)(MULT_SIZE-1) & MULT_33(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(53)(MULT_SIZE-1) & MULT_34(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(54)<=signed(MULT_33(54)(MULT_SIZE-1) & MULT_33(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(54)(MULT_SIZE-1) & MULT_34(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(55)<=signed(MULT_33(55)(MULT_SIZE-1) & MULT_33(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(55)(MULT_SIZE-1) & MULT_34(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(56)<=signed(MULT_33(56)(MULT_SIZE-1) & MULT_33(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(56)(MULT_SIZE-1) & MULT_34(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(57)<=signed(MULT_33(57)(MULT_SIZE-1) & MULT_33(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(57)(MULT_SIZE-1) & MULT_34(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(58)<=signed(MULT_33(58)(MULT_SIZE-1) & MULT_33(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(58)(MULT_SIZE-1) & MULT_34(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(59)<=signed(MULT_33(59)(MULT_SIZE-1) & MULT_33(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(59)(MULT_SIZE-1) & MULT_34(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(60)<=signed(MULT_33(60)(MULT_SIZE-1) & MULT_33(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(60)(MULT_SIZE-1) & MULT_34(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(61)<=signed(MULT_33(61)(MULT_SIZE-1) & MULT_33(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(61)(MULT_SIZE-1) & MULT_34(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(62)<=signed(MULT_33(62)(MULT_SIZE-1) & MULT_33(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(62)(MULT_SIZE-1) & MULT_34(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(63)<=signed(MULT_33(63)(MULT_SIZE-1) & MULT_33(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(63)(MULT_SIZE-1) & MULT_34(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(64)<=signed(MULT_33(64)(MULT_SIZE-1) & MULT_33(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(64)(MULT_SIZE-1) & MULT_34(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(65)<=signed(MULT_33(65)(MULT_SIZE-1) & MULT_33(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(65)(MULT_SIZE-1) & MULT_34(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(66)<=signed(MULT_33(66)(MULT_SIZE-1) & MULT_33(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(66)(MULT_SIZE-1) & MULT_34(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(67)<=signed(MULT_33(67)(MULT_SIZE-1) & MULT_33(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(67)(MULT_SIZE-1) & MULT_34(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(68)<=signed(MULT_33(68)(MULT_SIZE-1) & MULT_33(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(68)(MULT_SIZE-1) & MULT_34(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(69)<=signed(MULT_33(69)(MULT_SIZE-1) & MULT_33(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(69)(MULT_SIZE-1) & MULT_34(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(70)<=signed(MULT_33(70)(MULT_SIZE-1) & MULT_33(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(70)(MULT_SIZE-1) & MULT_34(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(71)<=signed(MULT_33(71)(MULT_SIZE-1) & MULT_33(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(71)(MULT_SIZE-1) & MULT_34(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(72)<=signed(MULT_33(72)(MULT_SIZE-1) & MULT_33(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(72)(MULT_SIZE-1) & MULT_34(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(73)<=signed(MULT_33(73)(MULT_SIZE-1) & MULT_33(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(73)(MULT_SIZE-1) & MULT_34(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(74)<=signed(MULT_33(74)(MULT_SIZE-1) & MULT_33(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(74)(MULT_SIZE-1) & MULT_34(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(75)<=signed(MULT_33(75)(MULT_SIZE-1) & MULT_33(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(75)(MULT_SIZE-1) & MULT_34(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(76)<=signed(MULT_33(76)(MULT_SIZE-1) & MULT_33(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(76)(MULT_SIZE-1) & MULT_34(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(77)<=signed(MULT_33(77)(MULT_SIZE-1) & MULT_33(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(77)(MULT_SIZE-1) & MULT_34(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(78)<=signed(MULT_33(78)(MULT_SIZE-1) & MULT_33(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(78)(MULT_SIZE-1) & MULT_34(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(79)<=signed(MULT_33(79)(MULT_SIZE-1) & MULT_33(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(79)(MULT_SIZE-1) & MULT_34(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(80)<=signed(MULT_33(80)(MULT_SIZE-1) & MULT_33(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(80)(MULT_SIZE-1) & MULT_34(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(81)<=signed(MULT_33(81)(MULT_SIZE-1) & MULT_33(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(81)(MULT_SIZE-1) & MULT_34(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(82)<=signed(MULT_33(82)(MULT_SIZE-1) & MULT_33(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(82)(MULT_SIZE-1) & MULT_34(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_17(83)<=signed(MULT_33(83)(MULT_SIZE-1) & MULT_33(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_34(83)(MULT_SIZE-1) & MULT_34(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_18(0)<=signed(MULT_35(0)(MULT_SIZE-1) & MULT_35(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(0)(MULT_SIZE-1) & MULT_36(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(1)<=signed(MULT_35(1)(MULT_SIZE-1) & MULT_35(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(1)(MULT_SIZE-1) & MULT_36(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(2)<=signed(MULT_35(2)(MULT_SIZE-1) & MULT_35(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(2)(MULT_SIZE-1) & MULT_36(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(3)<=signed(MULT_35(3)(MULT_SIZE-1) & MULT_35(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(3)(MULT_SIZE-1) & MULT_36(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(4)<=signed(MULT_35(4)(MULT_SIZE-1) & MULT_35(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(4)(MULT_SIZE-1) & MULT_36(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(5)<=signed(MULT_35(5)(MULT_SIZE-1) & MULT_35(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(5)(MULT_SIZE-1) & MULT_36(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(6)<=signed(MULT_35(6)(MULT_SIZE-1) & MULT_35(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(6)(MULT_SIZE-1) & MULT_36(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(7)<=signed(MULT_35(7)(MULT_SIZE-1) & MULT_35(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(7)(MULT_SIZE-1) & MULT_36(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(8)<=signed(MULT_35(8)(MULT_SIZE-1) & MULT_35(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(8)(MULT_SIZE-1) & MULT_36(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(9)<=signed(MULT_35(9)(MULT_SIZE-1) & MULT_35(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(9)(MULT_SIZE-1) & MULT_36(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(10)<=signed(MULT_35(10)(MULT_SIZE-1) & MULT_35(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(10)(MULT_SIZE-1) & MULT_36(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(11)<=signed(MULT_35(11)(MULT_SIZE-1) & MULT_35(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(11)(MULT_SIZE-1) & MULT_36(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(12)<=signed(MULT_35(12)(MULT_SIZE-1) & MULT_35(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(12)(MULT_SIZE-1) & MULT_36(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(13)<=signed(MULT_35(13)(MULT_SIZE-1) & MULT_35(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(13)(MULT_SIZE-1) & MULT_36(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(14)<=signed(MULT_35(14)(MULT_SIZE-1) & MULT_35(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(14)(MULT_SIZE-1) & MULT_36(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(15)<=signed(MULT_35(15)(MULT_SIZE-1) & MULT_35(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(15)(MULT_SIZE-1) & MULT_36(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(16)<=signed(MULT_35(16)(MULT_SIZE-1) & MULT_35(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(16)(MULT_SIZE-1) & MULT_36(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(17)<=signed(MULT_35(17)(MULT_SIZE-1) & MULT_35(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(17)(MULT_SIZE-1) & MULT_36(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(18)<=signed(MULT_35(18)(MULT_SIZE-1) & MULT_35(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(18)(MULT_SIZE-1) & MULT_36(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(19)<=signed(MULT_35(19)(MULT_SIZE-1) & MULT_35(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(19)(MULT_SIZE-1) & MULT_36(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(20)<=signed(MULT_35(20)(MULT_SIZE-1) & MULT_35(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(20)(MULT_SIZE-1) & MULT_36(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(21)<=signed(MULT_35(21)(MULT_SIZE-1) & MULT_35(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(21)(MULT_SIZE-1) & MULT_36(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(22)<=signed(MULT_35(22)(MULT_SIZE-1) & MULT_35(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(22)(MULT_SIZE-1) & MULT_36(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(23)<=signed(MULT_35(23)(MULT_SIZE-1) & MULT_35(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(23)(MULT_SIZE-1) & MULT_36(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(24)<=signed(MULT_35(24)(MULT_SIZE-1) & MULT_35(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(24)(MULT_SIZE-1) & MULT_36(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(25)<=signed(MULT_35(25)(MULT_SIZE-1) & MULT_35(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(25)(MULT_SIZE-1) & MULT_36(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(26)<=signed(MULT_35(26)(MULT_SIZE-1) & MULT_35(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(26)(MULT_SIZE-1) & MULT_36(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(27)<=signed(MULT_35(27)(MULT_SIZE-1) & MULT_35(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(27)(MULT_SIZE-1) & MULT_36(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(28)<=signed(MULT_35(28)(MULT_SIZE-1) & MULT_35(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(28)(MULT_SIZE-1) & MULT_36(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(29)<=signed(MULT_35(29)(MULT_SIZE-1) & MULT_35(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(29)(MULT_SIZE-1) & MULT_36(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(30)<=signed(MULT_35(30)(MULT_SIZE-1) & MULT_35(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(30)(MULT_SIZE-1) & MULT_36(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(31)<=signed(MULT_35(31)(MULT_SIZE-1) & MULT_35(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(31)(MULT_SIZE-1) & MULT_36(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(32)<=signed(MULT_35(32)(MULT_SIZE-1) & MULT_35(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(32)(MULT_SIZE-1) & MULT_36(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(33)<=signed(MULT_35(33)(MULT_SIZE-1) & MULT_35(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(33)(MULT_SIZE-1) & MULT_36(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(34)<=signed(MULT_35(34)(MULT_SIZE-1) & MULT_35(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(34)(MULT_SIZE-1) & MULT_36(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(35)<=signed(MULT_35(35)(MULT_SIZE-1) & MULT_35(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(35)(MULT_SIZE-1) & MULT_36(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(36)<=signed(MULT_35(36)(MULT_SIZE-1) & MULT_35(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(36)(MULT_SIZE-1) & MULT_36(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(37)<=signed(MULT_35(37)(MULT_SIZE-1) & MULT_35(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(37)(MULT_SIZE-1) & MULT_36(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(38)<=signed(MULT_35(38)(MULT_SIZE-1) & MULT_35(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(38)(MULT_SIZE-1) & MULT_36(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(39)<=signed(MULT_35(39)(MULT_SIZE-1) & MULT_35(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(39)(MULT_SIZE-1) & MULT_36(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(40)<=signed(MULT_35(40)(MULT_SIZE-1) & MULT_35(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(40)(MULT_SIZE-1) & MULT_36(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(41)<=signed(MULT_35(41)(MULT_SIZE-1) & MULT_35(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(41)(MULT_SIZE-1) & MULT_36(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(42)<=signed(MULT_35(42)(MULT_SIZE-1) & MULT_35(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(42)(MULT_SIZE-1) & MULT_36(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(43)<=signed(MULT_35(43)(MULT_SIZE-1) & MULT_35(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(43)(MULT_SIZE-1) & MULT_36(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(44)<=signed(MULT_35(44)(MULT_SIZE-1) & MULT_35(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(44)(MULT_SIZE-1) & MULT_36(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(45)<=signed(MULT_35(45)(MULT_SIZE-1) & MULT_35(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(45)(MULT_SIZE-1) & MULT_36(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(46)<=signed(MULT_35(46)(MULT_SIZE-1) & MULT_35(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(46)(MULT_SIZE-1) & MULT_36(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(47)<=signed(MULT_35(47)(MULT_SIZE-1) & MULT_35(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(47)(MULT_SIZE-1) & MULT_36(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(48)<=signed(MULT_35(48)(MULT_SIZE-1) & MULT_35(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(48)(MULT_SIZE-1) & MULT_36(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(49)<=signed(MULT_35(49)(MULT_SIZE-1) & MULT_35(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(49)(MULT_SIZE-1) & MULT_36(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(50)<=signed(MULT_35(50)(MULT_SIZE-1) & MULT_35(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(50)(MULT_SIZE-1) & MULT_36(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(51)<=signed(MULT_35(51)(MULT_SIZE-1) & MULT_35(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(51)(MULT_SIZE-1) & MULT_36(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(52)<=signed(MULT_35(52)(MULT_SIZE-1) & MULT_35(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(52)(MULT_SIZE-1) & MULT_36(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(53)<=signed(MULT_35(53)(MULT_SIZE-1) & MULT_35(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(53)(MULT_SIZE-1) & MULT_36(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(54)<=signed(MULT_35(54)(MULT_SIZE-1) & MULT_35(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(54)(MULT_SIZE-1) & MULT_36(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(55)<=signed(MULT_35(55)(MULT_SIZE-1) & MULT_35(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(55)(MULT_SIZE-1) & MULT_36(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(56)<=signed(MULT_35(56)(MULT_SIZE-1) & MULT_35(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(56)(MULT_SIZE-1) & MULT_36(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(57)<=signed(MULT_35(57)(MULT_SIZE-1) & MULT_35(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(57)(MULT_SIZE-1) & MULT_36(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(58)<=signed(MULT_35(58)(MULT_SIZE-1) & MULT_35(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(58)(MULT_SIZE-1) & MULT_36(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(59)<=signed(MULT_35(59)(MULT_SIZE-1) & MULT_35(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(59)(MULT_SIZE-1) & MULT_36(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(60)<=signed(MULT_35(60)(MULT_SIZE-1) & MULT_35(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(60)(MULT_SIZE-1) & MULT_36(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(61)<=signed(MULT_35(61)(MULT_SIZE-1) & MULT_35(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(61)(MULT_SIZE-1) & MULT_36(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(62)<=signed(MULT_35(62)(MULT_SIZE-1) & MULT_35(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(62)(MULT_SIZE-1) & MULT_36(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(63)<=signed(MULT_35(63)(MULT_SIZE-1) & MULT_35(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(63)(MULT_SIZE-1) & MULT_36(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(64)<=signed(MULT_35(64)(MULT_SIZE-1) & MULT_35(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(64)(MULT_SIZE-1) & MULT_36(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(65)<=signed(MULT_35(65)(MULT_SIZE-1) & MULT_35(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(65)(MULT_SIZE-1) & MULT_36(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(66)<=signed(MULT_35(66)(MULT_SIZE-1) & MULT_35(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(66)(MULT_SIZE-1) & MULT_36(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(67)<=signed(MULT_35(67)(MULT_SIZE-1) & MULT_35(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(67)(MULT_SIZE-1) & MULT_36(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(68)<=signed(MULT_35(68)(MULT_SIZE-1) & MULT_35(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(68)(MULT_SIZE-1) & MULT_36(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(69)<=signed(MULT_35(69)(MULT_SIZE-1) & MULT_35(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(69)(MULT_SIZE-1) & MULT_36(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(70)<=signed(MULT_35(70)(MULT_SIZE-1) & MULT_35(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(70)(MULT_SIZE-1) & MULT_36(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(71)<=signed(MULT_35(71)(MULT_SIZE-1) & MULT_35(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(71)(MULT_SIZE-1) & MULT_36(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(72)<=signed(MULT_35(72)(MULT_SIZE-1) & MULT_35(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(72)(MULT_SIZE-1) & MULT_36(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(73)<=signed(MULT_35(73)(MULT_SIZE-1) & MULT_35(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(73)(MULT_SIZE-1) & MULT_36(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(74)<=signed(MULT_35(74)(MULT_SIZE-1) & MULT_35(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(74)(MULT_SIZE-1) & MULT_36(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(75)<=signed(MULT_35(75)(MULT_SIZE-1) & MULT_35(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(75)(MULT_SIZE-1) & MULT_36(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(76)<=signed(MULT_35(76)(MULT_SIZE-1) & MULT_35(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(76)(MULT_SIZE-1) & MULT_36(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(77)<=signed(MULT_35(77)(MULT_SIZE-1) & MULT_35(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(77)(MULT_SIZE-1) & MULT_36(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(78)<=signed(MULT_35(78)(MULT_SIZE-1) & MULT_35(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(78)(MULT_SIZE-1) & MULT_36(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(79)<=signed(MULT_35(79)(MULT_SIZE-1) & MULT_35(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(79)(MULT_SIZE-1) & MULT_36(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(80)<=signed(MULT_35(80)(MULT_SIZE-1) & MULT_35(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(80)(MULT_SIZE-1) & MULT_36(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(81)<=signed(MULT_35(81)(MULT_SIZE-1) & MULT_35(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(81)(MULT_SIZE-1) & MULT_36(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(82)<=signed(MULT_35(82)(MULT_SIZE-1) & MULT_35(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(82)(MULT_SIZE-1) & MULT_36(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_18(83)<=signed(MULT_35(83)(MULT_SIZE-1) & MULT_35(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_36(83)(MULT_SIZE-1) & MULT_36(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_19(0)<=signed(MULT_37(0)(MULT_SIZE-1) & MULT_37(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(0)(MULT_SIZE-1) & MULT_38(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(1)<=signed(MULT_37(1)(MULT_SIZE-1) & MULT_37(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(1)(MULT_SIZE-1) & MULT_38(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(2)<=signed(MULT_37(2)(MULT_SIZE-1) & MULT_37(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(2)(MULT_SIZE-1) & MULT_38(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(3)<=signed(MULT_37(3)(MULT_SIZE-1) & MULT_37(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(3)(MULT_SIZE-1) & MULT_38(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(4)<=signed(MULT_37(4)(MULT_SIZE-1) & MULT_37(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(4)(MULT_SIZE-1) & MULT_38(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(5)<=signed(MULT_37(5)(MULT_SIZE-1) & MULT_37(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(5)(MULT_SIZE-1) & MULT_38(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(6)<=signed(MULT_37(6)(MULT_SIZE-1) & MULT_37(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(6)(MULT_SIZE-1) & MULT_38(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(7)<=signed(MULT_37(7)(MULT_SIZE-1) & MULT_37(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(7)(MULT_SIZE-1) & MULT_38(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(8)<=signed(MULT_37(8)(MULT_SIZE-1) & MULT_37(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(8)(MULT_SIZE-1) & MULT_38(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(9)<=signed(MULT_37(9)(MULT_SIZE-1) & MULT_37(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(9)(MULT_SIZE-1) & MULT_38(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(10)<=signed(MULT_37(10)(MULT_SIZE-1) & MULT_37(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(10)(MULT_SIZE-1) & MULT_38(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(11)<=signed(MULT_37(11)(MULT_SIZE-1) & MULT_37(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(11)(MULT_SIZE-1) & MULT_38(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(12)<=signed(MULT_37(12)(MULT_SIZE-1) & MULT_37(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(12)(MULT_SIZE-1) & MULT_38(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(13)<=signed(MULT_37(13)(MULT_SIZE-1) & MULT_37(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(13)(MULT_SIZE-1) & MULT_38(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(14)<=signed(MULT_37(14)(MULT_SIZE-1) & MULT_37(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(14)(MULT_SIZE-1) & MULT_38(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(15)<=signed(MULT_37(15)(MULT_SIZE-1) & MULT_37(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(15)(MULT_SIZE-1) & MULT_38(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(16)<=signed(MULT_37(16)(MULT_SIZE-1) & MULT_37(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(16)(MULT_SIZE-1) & MULT_38(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(17)<=signed(MULT_37(17)(MULT_SIZE-1) & MULT_37(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(17)(MULT_SIZE-1) & MULT_38(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(18)<=signed(MULT_37(18)(MULT_SIZE-1) & MULT_37(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(18)(MULT_SIZE-1) & MULT_38(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(19)<=signed(MULT_37(19)(MULT_SIZE-1) & MULT_37(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(19)(MULT_SIZE-1) & MULT_38(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(20)<=signed(MULT_37(20)(MULT_SIZE-1) & MULT_37(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(20)(MULT_SIZE-1) & MULT_38(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(21)<=signed(MULT_37(21)(MULT_SIZE-1) & MULT_37(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(21)(MULT_SIZE-1) & MULT_38(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(22)<=signed(MULT_37(22)(MULT_SIZE-1) & MULT_37(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(22)(MULT_SIZE-1) & MULT_38(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(23)<=signed(MULT_37(23)(MULT_SIZE-1) & MULT_37(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(23)(MULT_SIZE-1) & MULT_38(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(24)<=signed(MULT_37(24)(MULT_SIZE-1) & MULT_37(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(24)(MULT_SIZE-1) & MULT_38(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(25)<=signed(MULT_37(25)(MULT_SIZE-1) & MULT_37(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(25)(MULT_SIZE-1) & MULT_38(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(26)<=signed(MULT_37(26)(MULT_SIZE-1) & MULT_37(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(26)(MULT_SIZE-1) & MULT_38(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(27)<=signed(MULT_37(27)(MULT_SIZE-1) & MULT_37(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(27)(MULT_SIZE-1) & MULT_38(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(28)<=signed(MULT_37(28)(MULT_SIZE-1) & MULT_37(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(28)(MULT_SIZE-1) & MULT_38(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(29)<=signed(MULT_37(29)(MULT_SIZE-1) & MULT_37(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(29)(MULT_SIZE-1) & MULT_38(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(30)<=signed(MULT_37(30)(MULT_SIZE-1) & MULT_37(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(30)(MULT_SIZE-1) & MULT_38(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(31)<=signed(MULT_37(31)(MULT_SIZE-1) & MULT_37(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(31)(MULT_SIZE-1) & MULT_38(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(32)<=signed(MULT_37(32)(MULT_SIZE-1) & MULT_37(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(32)(MULT_SIZE-1) & MULT_38(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(33)<=signed(MULT_37(33)(MULT_SIZE-1) & MULT_37(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(33)(MULT_SIZE-1) & MULT_38(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(34)<=signed(MULT_37(34)(MULT_SIZE-1) & MULT_37(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(34)(MULT_SIZE-1) & MULT_38(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(35)<=signed(MULT_37(35)(MULT_SIZE-1) & MULT_37(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(35)(MULT_SIZE-1) & MULT_38(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(36)<=signed(MULT_37(36)(MULT_SIZE-1) & MULT_37(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(36)(MULT_SIZE-1) & MULT_38(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(37)<=signed(MULT_37(37)(MULT_SIZE-1) & MULT_37(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(37)(MULT_SIZE-1) & MULT_38(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(38)<=signed(MULT_37(38)(MULT_SIZE-1) & MULT_37(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(38)(MULT_SIZE-1) & MULT_38(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(39)<=signed(MULT_37(39)(MULT_SIZE-1) & MULT_37(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(39)(MULT_SIZE-1) & MULT_38(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(40)<=signed(MULT_37(40)(MULT_SIZE-1) & MULT_37(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(40)(MULT_SIZE-1) & MULT_38(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(41)<=signed(MULT_37(41)(MULT_SIZE-1) & MULT_37(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(41)(MULT_SIZE-1) & MULT_38(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(42)<=signed(MULT_37(42)(MULT_SIZE-1) & MULT_37(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(42)(MULT_SIZE-1) & MULT_38(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(43)<=signed(MULT_37(43)(MULT_SIZE-1) & MULT_37(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(43)(MULT_SIZE-1) & MULT_38(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(44)<=signed(MULT_37(44)(MULT_SIZE-1) & MULT_37(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(44)(MULT_SIZE-1) & MULT_38(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(45)<=signed(MULT_37(45)(MULT_SIZE-1) & MULT_37(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(45)(MULT_SIZE-1) & MULT_38(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(46)<=signed(MULT_37(46)(MULT_SIZE-1) & MULT_37(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(46)(MULT_SIZE-1) & MULT_38(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(47)<=signed(MULT_37(47)(MULT_SIZE-1) & MULT_37(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(47)(MULT_SIZE-1) & MULT_38(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(48)<=signed(MULT_37(48)(MULT_SIZE-1) & MULT_37(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(48)(MULT_SIZE-1) & MULT_38(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(49)<=signed(MULT_37(49)(MULT_SIZE-1) & MULT_37(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(49)(MULT_SIZE-1) & MULT_38(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(50)<=signed(MULT_37(50)(MULT_SIZE-1) & MULT_37(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(50)(MULT_SIZE-1) & MULT_38(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(51)<=signed(MULT_37(51)(MULT_SIZE-1) & MULT_37(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(51)(MULT_SIZE-1) & MULT_38(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(52)<=signed(MULT_37(52)(MULT_SIZE-1) & MULT_37(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(52)(MULT_SIZE-1) & MULT_38(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(53)<=signed(MULT_37(53)(MULT_SIZE-1) & MULT_37(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(53)(MULT_SIZE-1) & MULT_38(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(54)<=signed(MULT_37(54)(MULT_SIZE-1) & MULT_37(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(54)(MULT_SIZE-1) & MULT_38(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(55)<=signed(MULT_37(55)(MULT_SIZE-1) & MULT_37(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(55)(MULT_SIZE-1) & MULT_38(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(56)<=signed(MULT_37(56)(MULT_SIZE-1) & MULT_37(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(56)(MULT_SIZE-1) & MULT_38(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(57)<=signed(MULT_37(57)(MULT_SIZE-1) & MULT_37(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(57)(MULT_SIZE-1) & MULT_38(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(58)<=signed(MULT_37(58)(MULT_SIZE-1) & MULT_37(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(58)(MULT_SIZE-1) & MULT_38(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(59)<=signed(MULT_37(59)(MULT_SIZE-1) & MULT_37(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(59)(MULT_SIZE-1) & MULT_38(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(60)<=signed(MULT_37(60)(MULT_SIZE-1) & MULT_37(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(60)(MULT_SIZE-1) & MULT_38(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(61)<=signed(MULT_37(61)(MULT_SIZE-1) & MULT_37(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(61)(MULT_SIZE-1) & MULT_38(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(62)<=signed(MULT_37(62)(MULT_SIZE-1) & MULT_37(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(62)(MULT_SIZE-1) & MULT_38(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(63)<=signed(MULT_37(63)(MULT_SIZE-1) & MULT_37(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(63)(MULT_SIZE-1) & MULT_38(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(64)<=signed(MULT_37(64)(MULT_SIZE-1) & MULT_37(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(64)(MULT_SIZE-1) & MULT_38(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(65)<=signed(MULT_37(65)(MULT_SIZE-1) & MULT_37(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(65)(MULT_SIZE-1) & MULT_38(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(66)<=signed(MULT_37(66)(MULT_SIZE-1) & MULT_37(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(66)(MULT_SIZE-1) & MULT_38(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(67)<=signed(MULT_37(67)(MULT_SIZE-1) & MULT_37(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(67)(MULT_SIZE-1) & MULT_38(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(68)<=signed(MULT_37(68)(MULT_SIZE-1) & MULT_37(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(68)(MULT_SIZE-1) & MULT_38(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(69)<=signed(MULT_37(69)(MULT_SIZE-1) & MULT_37(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(69)(MULT_SIZE-1) & MULT_38(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(70)<=signed(MULT_37(70)(MULT_SIZE-1) & MULT_37(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(70)(MULT_SIZE-1) & MULT_38(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(71)<=signed(MULT_37(71)(MULT_SIZE-1) & MULT_37(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(71)(MULT_SIZE-1) & MULT_38(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(72)<=signed(MULT_37(72)(MULT_SIZE-1) & MULT_37(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(72)(MULT_SIZE-1) & MULT_38(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(73)<=signed(MULT_37(73)(MULT_SIZE-1) & MULT_37(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(73)(MULT_SIZE-1) & MULT_38(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(74)<=signed(MULT_37(74)(MULT_SIZE-1) & MULT_37(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(74)(MULT_SIZE-1) & MULT_38(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(75)<=signed(MULT_37(75)(MULT_SIZE-1) & MULT_37(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(75)(MULT_SIZE-1) & MULT_38(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(76)<=signed(MULT_37(76)(MULT_SIZE-1) & MULT_37(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(76)(MULT_SIZE-1) & MULT_38(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(77)<=signed(MULT_37(77)(MULT_SIZE-1) & MULT_37(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(77)(MULT_SIZE-1) & MULT_38(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(78)<=signed(MULT_37(78)(MULT_SIZE-1) & MULT_37(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(78)(MULT_SIZE-1) & MULT_38(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(79)<=signed(MULT_37(79)(MULT_SIZE-1) & MULT_37(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(79)(MULT_SIZE-1) & MULT_38(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(80)<=signed(MULT_37(80)(MULT_SIZE-1) & MULT_37(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(80)(MULT_SIZE-1) & MULT_38(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(81)<=signed(MULT_37(81)(MULT_SIZE-1) & MULT_37(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(81)(MULT_SIZE-1) & MULT_38(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(82)<=signed(MULT_37(82)(MULT_SIZE-1) & MULT_37(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(82)(MULT_SIZE-1) & MULT_38(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_19(83)<=signed(MULT_37(83)(MULT_SIZE-1) & MULT_37(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_38(83)(MULT_SIZE-1) & MULT_38(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_20(0)<=signed(MULT_39(0)(MULT_SIZE-1) & MULT_39(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(0)(MULT_SIZE-1) & MULT_40(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(1)<=signed(MULT_39(1)(MULT_SIZE-1) & MULT_39(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(1)(MULT_SIZE-1) & MULT_40(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(2)<=signed(MULT_39(2)(MULT_SIZE-1) & MULT_39(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(2)(MULT_SIZE-1) & MULT_40(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(3)<=signed(MULT_39(3)(MULT_SIZE-1) & MULT_39(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(3)(MULT_SIZE-1) & MULT_40(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(4)<=signed(MULT_39(4)(MULT_SIZE-1) & MULT_39(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(4)(MULT_SIZE-1) & MULT_40(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(5)<=signed(MULT_39(5)(MULT_SIZE-1) & MULT_39(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(5)(MULT_SIZE-1) & MULT_40(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(6)<=signed(MULT_39(6)(MULT_SIZE-1) & MULT_39(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(6)(MULT_SIZE-1) & MULT_40(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(7)<=signed(MULT_39(7)(MULT_SIZE-1) & MULT_39(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(7)(MULT_SIZE-1) & MULT_40(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(8)<=signed(MULT_39(8)(MULT_SIZE-1) & MULT_39(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(8)(MULT_SIZE-1) & MULT_40(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(9)<=signed(MULT_39(9)(MULT_SIZE-1) & MULT_39(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(9)(MULT_SIZE-1) & MULT_40(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(10)<=signed(MULT_39(10)(MULT_SIZE-1) & MULT_39(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(10)(MULT_SIZE-1) & MULT_40(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(11)<=signed(MULT_39(11)(MULT_SIZE-1) & MULT_39(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(11)(MULT_SIZE-1) & MULT_40(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(12)<=signed(MULT_39(12)(MULT_SIZE-1) & MULT_39(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(12)(MULT_SIZE-1) & MULT_40(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(13)<=signed(MULT_39(13)(MULT_SIZE-1) & MULT_39(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(13)(MULT_SIZE-1) & MULT_40(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(14)<=signed(MULT_39(14)(MULT_SIZE-1) & MULT_39(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(14)(MULT_SIZE-1) & MULT_40(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(15)<=signed(MULT_39(15)(MULT_SIZE-1) & MULT_39(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(15)(MULT_SIZE-1) & MULT_40(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(16)<=signed(MULT_39(16)(MULT_SIZE-1) & MULT_39(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(16)(MULT_SIZE-1) & MULT_40(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(17)<=signed(MULT_39(17)(MULT_SIZE-1) & MULT_39(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(17)(MULT_SIZE-1) & MULT_40(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(18)<=signed(MULT_39(18)(MULT_SIZE-1) & MULT_39(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(18)(MULT_SIZE-1) & MULT_40(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(19)<=signed(MULT_39(19)(MULT_SIZE-1) & MULT_39(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(19)(MULT_SIZE-1) & MULT_40(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(20)<=signed(MULT_39(20)(MULT_SIZE-1) & MULT_39(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(20)(MULT_SIZE-1) & MULT_40(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(21)<=signed(MULT_39(21)(MULT_SIZE-1) & MULT_39(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(21)(MULT_SIZE-1) & MULT_40(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(22)<=signed(MULT_39(22)(MULT_SIZE-1) & MULT_39(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(22)(MULT_SIZE-1) & MULT_40(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(23)<=signed(MULT_39(23)(MULT_SIZE-1) & MULT_39(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(23)(MULT_SIZE-1) & MULT_40(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(24)<=signed(MULT_39(24)(MULT_SIZE-1) & MULT_39(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(24)(MULT_SIZE-1) & MULT_40(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(25)<=signed(MULT_39(25)(MULT_SIZE-1) & MULT_39(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(25)(MULT_SIZE-1) & MULT_40(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(26)<=signed(MULT_39(26)(MULT_SIZE-1) & MULT_39(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(26)(MULT_SIZE-1) & MULT_40(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(27)<=signed(MULT_39(27)(MULT_SIZE-1) & MULT_39(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(27)(MULT_SIZE-1) & MULT_40(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(28)<=signed(MULT_39(28)(MULT_SIZE-1) & MULT_39(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(28)(MULT_SIZE-1) & MULT_40(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(29)<=signed(MULT_39(29)(MULT_SIZE-1) & MULT_39(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(29)(MULT_SIZE-1) & MULT_40(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(30)<=signed(MULT_39(30)(MULT_SIZE-1) & MULT_39(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(30)(MULT_SIZE-1) & MULT_40(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(31)<=signed(MULT_39(31)(MULT_SIZE-1) & MULT_39(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(31)(MULT_SIZE-1) & MULT_40(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(32)<=signed(MULT_39(32)(MULT_SIZE-1) & MULT_39(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(32)(MULT_SIZE-1) & MULT_40(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(33)<=signed(MULT_39(33)(MULT_SIZE-1) & MULT_39(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(33)(MULT_SIZE-1) & MULT_40(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(34)<=signed(MULT_39(34)(MULT_SIZE-1) & MULT_39(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(34)(MULT_SIZE-1) & MULT_40(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(35)<=signed(MULT_39(35)(MULT_SIZE-1) & MULT_39(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(35)(MULT_SIZE-1) & MULT_40(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(36)<=signed(MULT_39(36)(MULT_SIZE-1) & MULT_39(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(36)(MULT_SIZE-1) & MULT_40(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(37)<=signed(MULT_39(37)(MULT_SIZE-1) & MULT_39(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(37)(MULT_SIZE-1) & MULT_40(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(38)<=signed(MULT_39(38)(MULT_SIZE-1) & MULT_39(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(38)(MULT_SIZE-1) & MULT_40(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(39)<=signed(MULT_39(39)(MULT_SIZE-1) & MULT_39(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(39)(MULT_SIZE-1) & MULT_40(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(40)<=signed(MULT_39(40)(MULT_SIZE-1) & MULT_39(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(40)(MULT_SIZE-1) & MULT_40(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(41)<=signed(MULT_39(41)(MULT_SIZE-1) & MULT_39(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(41)(MULT_SIZE-1) & MULT_40(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(42)<=signed(MULT_39(42)(MULT_SIZE-1) & MULT_39(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(42)(MULT_SIZE-1) & MULT_40(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(43)<=signed(MULT_39(43)(MULT_SIZE-1) & MULT_39(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(43)(MULT_SIZE-1) & MULT_40(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(44)<=signed(MULT_39(44)(MULT_SIZE-1) & MULT_39(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(44)(MULT_SIZE-1) & MULT_40(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(45)<=signed(MULT_39(45)(MULT_SIZE-1) & MULT_39(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(45)(MULT_SIZE-1) & MULT_40(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(46)<=signed(MULT_39(46)(MULT_SIZE-1) & MULT_39(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(46)(MULT_SIZE-1) & MULT_40(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(47)<=signed(MULT_39(47)(MULT_SIZE-1) & MULT_39(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(47)(MULT_SIZE-1) & MULT_40(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(48)<=signed(MULT_39(48)(MULT_SIZE-1) & MULT_39(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(48)(MULT_SIZE-1) & MULT_40(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(49)<=signed(MULT_39(49)(MULT_SIZE-1) & MULT_39(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(49)(MULT_SIZE-1) & MULT_40(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(50)<=signed(MULT_39(50)(MULT_SIZE-1) & MULT_39(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(50)(MULT_SIZE-1) & MULT_40(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(51)<=signed(MULT_39(51)(MULT_SIZE-1) & MULT_39(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(51)(MULT_SIZE-1) & MULT_40(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(52)<=signed(MULT_39(52)(MULT_SIZE-1) & MULT_39(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(52)(MULT_SIZE-1) & MULT_40(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(53)<=signed(MULT_39(53)(MULT_SIZE-1) & MULT_39(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(53)(MULT_SIZE-1) & MULT_40(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(54)<=signed(MULT_39(54)(MULT_SIZE-1) & MULT_39(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(54)(MULT_SIZE-1) & MULT_40(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(55)<=signed(MULT_39(55)(MULT_SIZE-1) & MULT_39(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(55)(MULT_SIZE-1) & MULT_40(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(56)<=signed(MULT_39(56)(MULT_SIZE-1) & MULT_39(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(56)(MULT_SIZE-1) & MULT_40(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(57)<=signed(MULT_39(57)(MULT_SIZE-1) & MULT_39(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(57)(MULT_SIZE-1) & MULT_40(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(58)<=signed(MULT_39(58)(MULT_SIZE-1) & MULT_39(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(58)(MULT_SIZE-1) & MULT_40(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(59)<=signed(MULT_39(59)(MULT_SIZE-1) & MULT_39(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(59)(MULT_SIZE-1) & MULT_40(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(60)<=signed(MULT_39(60)(MULT_SIZE-1) & MULT_39(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(60)(MULT_SIZE-1) & MULT_40(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(61)<=signed(MULT_39(61)(MULT_SIZE-1) & MULT_39(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(61)(MULT_SIZE-1) & MULT_40(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(62)<=signed(MULT_39(62)(MULT_SIZE-1) & MULT_39(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(62)(MULT_SIZE-1) & MULT_40(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(63)<=signed(MULT_39(63)(MULT_SIZE-1) & MULT_39(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(63)(MULT_SIZE-1) & MULT_40(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(64)<=signed(MULT_39(64)(MULT_SIZE-1) & MULT_39(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(64)(MULT_SIZE-1) & MULT_40(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(65)<=signed(MULT_39(65)(MULT_SIZE-1) & MULT_39(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(65)(MULT_SIZE-1) & MULT_40(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(66)<=signed(MULT_39(66)(MULT_SIZE-1) & MULT_39(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(66)(MULT_SIZE-1) & MULT_40(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(67)<=signed(MULT_39(67)(MULT_SIZE-1) & MULT_39(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(67)(MULT_SIZE-1) & MULT_40(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(68)<=signed(MULT_39(68)(MULT_SIZE-1) & MULT_39(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(68)(MULT_SIZE-1) & MULT_40(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(69)<=signed(MULT_39(69)(MULT_SIZE-1) & MULT_39(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(69)(MULT_SIZE-1) & MULT_40(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(70)<=signed(MULT_39(70)(MULT_SIZE-1) & MULT_39(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(70)(MULT_SIZE-1) & MULT_40(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(71)<=signed(MULT_39(71)(MULT_SIZE-1) & MULT_39(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(71)(MULT_SIZE-1) & MULT_40(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(72)<=signed(MULT_39(72)(MULT_SIZE-1) & MULT_39(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(72)(MULT_SIZE-1) & MULT_40(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(73)<=signed(MULT_39(73)(MULT_SIZE-1) & MULT_39(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(73)(MULT_SIZE-1) & MULT_40(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(74)<=signed(MULT_39(74)(MULT_SIZE-1) & MULT_39(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(74)(MULT_SIZE-1) & MULT_40(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(75)<=signed(MULT_39(75)(MULT_SIZE-1) & MULT_39(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(75)(MULT_SIZE-1) & MULT_40(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(76)<=signed(MULT_39(76)(MULT_SIZE-1) & MULT_39(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(76)(MULT_SIZE-1) & MULT_40(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(77)<=signed(MULT_39(77)(MULT_SIZE-1) & MULT_39(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(77)(MULT_SIZE-1) & MULT_40(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(78)<=signed(MULT_39(78)(MULT_SIZE-1) & MULT_39(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(78)(MULT_SIZE-1) & MULT_40(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(79)<=signed(MULT_39(79)(MULT_SIZE-1) & MULT_39(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(79)(MULT_SIZE-1) & MULT_40(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(80)<=signed(MULT_39(80)(MULT_SIZE-1) & MULT_39(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(80)(MULT_SIZE-1) & MULT_40(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(81)<=signed(MULT_39(81)(MULT_SIZE-1) & MULT_39(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(81)(MULT_SIZE-1) & MULT_40(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(82)<=signed(MULT_39(82)(MULT_SIZE-1) & MULT_39(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(82)(MULT_SIZE-1) & MULT_40(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_20(83)<=signed(MULT_39(83)(MULT_SIZE-1) & MULT_39(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_40(83)(MULT_SIZE-1) & MULT_40(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_21(0)<=signed(MULT_41(0)(MULT_SIZE-1) & MULT_41(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(0)(MULT_SIZE-1) & MULT_42(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(1)<=signed(MULT_41(1)(MULT_SIZE-1) & MULT_41(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(1)(MULT_SIZE-1) & MULT_42(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(2)<=signed(MULT_41(2)(MULT_SIZE-1) & MULT_41(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(2)(MULT_SIZE-1) & MULT_42(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(3)<=signed(MULT_41(3)(MULT_SIZE-1) & MULT_41(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(3)(MULT_SIZE-1) & MULT_42(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(4)<=signed(MULT_41(4)(MULT_SIZE-1) & MULT_41(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(4)(MULT_SIZE-1) & MULT_42(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(5)<=signed(MULT_41(5)(MULT_SIZE-1) & MULT_41(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(5)(MULT_SIZE-1) & MULT_42(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(6)<=signed(MULT_41(6)(MULT_SIZE-1) & MULT_41(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(6)(MULT_SIZE-1) & MULT_42(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(7)<=signed(MULT_41(7)(MULT_SIZE-1) & MULT_41(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(7)(MULT_SIZE-1) & MULT_42(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(8)<=signed(MULT_41(8)(MULT_SIZE-1) & MULT_41(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(8)(MULT_SIZE-1) & MULT_42(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(9)<=signed(MULT_41(9)(MULT_SIZE-1) & MULT_41(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(9)(MULT_SIZE-1) & MULT_42(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(10)<=signed(MULT_41(10)(MULT_SIZE-1) & MULT_41(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(10)(MULT_SIZE-1) & MULT_42(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(11)<=signed(MULT_41(11)(MULT_SIZE-1) & MULT_41(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(11)(MULT_SIZE-1) & MULT_42(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(12)<=signed(MULT_41(12)(MULT_SIZE-1) & MULT_41(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(12)(MULT_SIZE-1) & MULT_42(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(13)<=signed(MULT_41(13)(MULT_SIZE-1) & MULT_41(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(13)(MULT_SIZE-1) & MULT_42(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(14)<=signed(MULT_41(14)(MULT_SIZE-1) & MULT_41(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(14)(MULT_SIZE-1) & MULT_42(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(15)<=signed(MULT_41(15)(MULT_SIZE-1) & MULT_41(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(15)(MULT_SIZE-1) & MULT_42(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(16)<=signed(MULT_41(16)(MULT_SIZE-1) & MULT_41(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(16)(MULT_SIZE-1) & MULT_42(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(17)<=signed(MULT_41(17)(MULT_SIZE-1) & MULT_41(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(17)(MULT_SIZE-1) & MULT_42(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(18)<=signed(MULT_41(18)(MULT_SIZE-1) & MULT_41(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(18)(MULT_SIZE-1) & MULT_42(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(19)<=signed(MULT_41(19)(MULT_SIZE-1) & MULT_41(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(19)(MULT_SIZE-1) & MULT_42(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(20)<=signed(MULT_41(20)(MULT_SIZE-1) & MULT_41(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(20)(MULT_SIZE-1) & MULT_42(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(21)<=signed(MULT_41(21)(MULT_SIZE-1) & MULT_41(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(21)(MULT_SIZE-1) & MULT_42(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(22)<=signed(MULT_41(22)(MULT_SIZE-1) & MULT_41(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(22)(MULT_SIZE-1) & MULT_42(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(23)<=signed(MULT_41(23)(MULT_SIZE-1) & MULT_41(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(23)(MULT_SIZE-1) & MULT_42(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(24)<=signed(MULT_41(24)(MULT_SIZE-1) & MULT_41(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(24)(MULT_SIZE-1) & MULT_42(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(25)<=signed(MULT_41(25)(MULT_SIZE-1) & MULT_41(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(25)(MULT_SIZE-1) & MULT_42(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(26)<=signed(MULT_41(26)(MULT_SIZE-1) & MULT_41(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(26)(MULT_SIZE-1) & MULT_42(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(27)<=signed(MULT_41(27)(MULT_SIZE-1) & MULT_41(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(27)(MULT_SIZE-1) & MULT_42(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(28)<=signed(MULT_41(28)(MULT_SIZE-1) & MULT_41(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(28)(MULT_SIZE-1) & MULT_42(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(29)<=signed(MULT_41(29)(MULT_SIZE-1) & MULT_41(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(29)(MULT_SIZE-1) & MULT_42(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(30)<=signed(MULT_41(30)(MULT_SIZE-1) & MULT_41(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(30)(MULT_SIZE-1) & MULT_42(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(31)<=signed(MULT_41(31)(MULT_SIZE-1) & MULT_41(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(31)(MULT_SIZE-1) & MULT_42(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(32)<=signed(MULT_41(32)(MULT_SIZE-1) & MULT_41(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(32)(MULT_SIZE-1) & MULT_42(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(33)<=signed(MULT_41(33)(MULT_SIZE-1) & MULT_41(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(33)(MULT_SIZE-1) & MULT_42(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(34)<=signed(MULT_41(34)(MULT_SIZE-1) & MULT_41(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(34)(MULT_SIZE-1) & MULT_42(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(35)<=signed(MULT_41(35)(MULT_SIZE-1) & MULT_41(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(35)(MULT_SIZE-1) & MULT_42(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(36)<=signed(MULT_41(36)(MULT_SIZE-1) & MULT_41(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(36)(MULT_SIZE-1) & MULT_42(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(37)<=signed(MULT_41(37)(MULT_SIZE-1) & MULT_41(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(37)(MULT_SIZE-1) & MULT_42(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(38)<=signed(MULT_41(38)(MULT_SIZE-1) & MULT_41(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(38)(MULT_SIZE-1) & MULT_42(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(39)<=signed(MULT_41(39)(MULT_SIZE-1) & MULT_41(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(39)(MULT_SIZE-1) & MULT_42(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(40)<=signed(MULT_41(40)(MULT_SIZE-1) & MULT_41(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(40)(MULT_SIZE-1) & MULT_42(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(41)<=signed(MULT_41(41)(MULT_SIZE-1) & MULT_41(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(41)(MULT_SIZE-1) & MULT_42(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(42)<=signed(MULT_41(42)(MULT_SIZE-1) & MULT_41(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(42)(MULT_SIZE-1) & MULT_42(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(43)<=signed(MULT_41(43)(MULT_SIZE-1) & MULT_41(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(43)(MULT_SIZE-1) & MULT_42(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(44)<=signed(MULT_41(44)(MULT_SIZE-1) & MULT_41(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(44)(MULT_SIZE-1) & MULT_42(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(45)<=signed(MULT_41(45)(MULT_SIZE-1) & MULT_41(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(45)(MULT_SIZE-1) & MULT_42(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(46)<=signed(MULT_41(46)(MULT_SIZE-1) & MULT_41(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(46)(MULT_SIZE-1) & MULT_42(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(47)<=signed(MULT_41(47)(MULT_SIZE-1) & MULT_41(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(47)(MULT_SIZE-1) & MULT_42(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(48)<=signed(MULT_41(48)(MULT_SIZE-1) & MULT_41(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(48)(MULT_SIZE-1) & MULT_42(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(49)<=signed(MULT_41(49)(MULT_SIZE-1) & MULT_41(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(49)(MULT_SIZE-1) & MULT_42(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(50)<=signed(MULT_41(50)(MULT_SIZE-1) & MULT_41(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(50)(MULT_SIZE-1) & MULT_42(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(51)<=signed(MULT_41(51)(MULT_SIZE-1) & MULT_41(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(51)(MULT_SIZE-1) & MULT_42(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(52)<=signed(MULT_41(52)(MULT_SIZE-1) & MULT_41(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(52)(MULT_SIZE-1) & MULT_42(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(53)<=signed(MULT_41(53)(MULT_SIZE-1) & MULT_41(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(53)(MULT_SIZE-1) & MULT_42(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(54)<=signed(MULT_41(54)(MULT_SIZE-1) & MULT_41(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(54)(MULT_SIZE-1) & MULT_42(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(55)<=signed(MULT_41(55)(MULT_SIZE-1) & MULT_41(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(55)(MULT_SIZE-1) & MULT_42(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(56)<=signed(MULT_41(56)(MULT_SIZE-1) & MULT_41(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(56)(MULT_SIZE-1) & MULT_42(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(57)<=signed(MULT_41(57)(MULT_SIZE-1) & MULT_41(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(57)(MULT_SIZE-1) & MULT_42(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(58)<=signed(MULT_41(58)(MULT_SIZE-1) & MULT_41(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(58)(MULT_SIZE-1) & MULT_42(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(59)<=signed(MULT_41(59)(MULT_SIZE-1) & MULT_41(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(59)(MULT_SIZE-1) & MULT_42(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(60)<=signed(MULT_41(60)(MULT_SIZE-1) & MULT_41(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(60)(MULT_SIZE-1) & MULT_42(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(61)<=signed(MULT_41(61)(MULT_SIZE-1) & MULT_41(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(61)(MULT_SIZE-1) & MULT_42(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(62)<=signed(MULT_41(62)(MULT_SIZE-1) & MULT_41(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(62)(MULT_SIZE-1) & MULT_42(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(63)<=signed(MULT_41(63)(MULT_SIZE-1) & MULT_41(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(63)(MULT_SIZE-1) & MULT_42(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(64)<=signed(MULT_41(64)(MULT_SIZE-1) & MULT_41(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(64)(MULT_SIZE-1) & MULT_42(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(65)<=signed(MULT_41(65)(MULT_SIZE-1) & MULT_41(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(65)(MULT_SIZE-1) & MULT_42(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(66)<=signed(MULT_41(66)(MULT_SIZE-1) & MULT_41(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(66)(MULT_SIZE-1) & MULT_42(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(67)<=signed(MULT_41(67)(MULT_SIZE-1) & MULT_41(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(67)(MULT_SIZE-1) & MULT_42(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(68)<=signed(MULT_41(68)(MULT_SIZE-1) & MULT_41(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(68)(MULT_SIZE-1) & MULT_42(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(69)<=signed(MULT_41(69)(MULT_SIZE-1) & MULT_41(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(69)(MULT_SIZE-1) & MULT_42(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(70)<=signed(MULT_41(70)(MULT_SIZE-1) & MULT_41(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(70)(MULT_SIZE-1) & MULT_42(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(71)<=signed(MULT_41(71)(MULT_SIZE-1) & MULT_41(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(71)(MULT_SIZE-1) & MULT_42(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(72)<=signed(MULT_41(72)(MULT_SIZE-1) & MULT_41(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(72)(MULT_SIZE-1) & MULT_42(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(73)<=signed(MULT_41(73)(MULT_SIZE-1) & MULT_41(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(73)(MULT_SIZE-1) & MULT_42(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(74)<=signed(MULT_41(74)(MULT_SIZE-1) & MULT_41(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(74)(MULT_SIZE-1) & MULT_42(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(75)<=signed(MULT_41(75)(MULT_SIZE-1) & MULT_41(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(75)(MULT_SIZE-1) & MULT_42(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(76)<=signed(MULT_41(76)(MULT_SIZE-1) & MULT_41(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(76)(MULT_SIZE-1) & MULT_42(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(77)<=signed(MULT_41(77)(MULT_SIZE-1) & MULT_41(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(77)(MULT_SIZE-1) & MULT_42(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(78)<=signed(MULT_41(78)(MULT_SIZE-1) & MULT_41(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(78)(MULT_SIZE-1) & MULT_42(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(79)<=signed(MULT_41(79)(MULT_SIZE-1) & MULT_41(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(79)(MULT_SIZE-1) & MULT_42(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(80)<=signed(MULT_41(80)(MULT_SIZE-1) & MULT_41(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(80)(MULT_SIZE-1) & MULT_42(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(81)<=signed(MULT_41(81)(MULT_SIZE-1) & MULT_41(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(81)(MULT_SIZE-1) & MULT_42(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(82)<=signed(MULT_41(82)(MULT_SIZE-1) & MULT_41(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(82)(MULT_SIZE-1) & MULT_42(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_21(83)<=signed(MULT_41(83)(MULT_SIZE-1) & MULT_41(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_42(83)(MULT_SIZE-1) & MULT_42(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_22(0)<=signed(MULT_43(0)(MULT_SIZE-1) & MULT_43(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(0)(MULT_SIZE-1) & MULT_44(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(1)<=signed(MULT_43(1)(MULT_SIZE-1) & MULT_43(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(1)(MULT_SIZE-1) & MULT_44(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(2)<=signed(MULT_43(2)(MULT_SIZE-1) & MULT_43(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(2)(MULT_SIZE-1) & MULT_44(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(3)<=signed(MULT_43(3)(MULT_SIZE-1) & MULT_43(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(3)(MULT_SIZE-1) & MULT_44(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(4)<=signed(MULT_43(4)(MULT_SIZE-1) & MULT_43(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(4)(MULT_SIZE-1) & MULT_44(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(5)<=signed(MULT_43(5)(MULT_SIZE-1) & MULT_43(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(5)(MULT_SIZE-1) & MULT_44(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(6)<=signed(MULT_43(6)(MULT_SIZE-1) & MULT_43(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(6)(MULT_SIZE-1) & MULT_44(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(7)<=signed(MULT_43(7)(MULT_SIZE-1) & MULT_43(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(7)(MULT_SIZE-1) & MULT_44(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(8)<=signed(MULT_43(8)(MULT_SIZE-1) & MULT_43(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(8)(MULT_SIZE-1) & MULT_44(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(9)<=signed(MULT_43(9)(MULT_SIZE-1) & MULT_43(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(9)(MULT_SIZE-1) & MULT_44(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(10)<=signed(MULT_43(10)(MULT_SIZE-1) & MULT_43(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(10)(MULT_SIZE-1) & MULT_44(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(11)<=signed(MULT_43(11)(MULT_SIZE-1) & MULT_43(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(11)(MULT_SIZE-1) & MULT_44(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(12)<=signed(MULT_43(12)(MULT_SIZE-1) & MULT_43(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(12)(MULT_SIZE-1) & MULT_44(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(13)<=signed(MULT_43(13)(MULT_SIZE-1) & MULT_43(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(13)(MULT_SIZE-1) & MULT_44(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(14)<=signed(MULT_43(14)(MULT_SIZE-1) & MULT_43(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(14)(MULT_SIZE-1) & MULT_44(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(15)<=signed(MULT_43(15)(MULT_SIZE-1) & MULT_43(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(15)(MULT_SIZE-1) & MULT_44(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(16)<=signed(MULT_43(16)(MULT_SIZE-1) & MULT_43(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(16)(MULT_SIZE-1) & MULT_44(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(17)<=signed(MULT_43(17)(MULT_SIZE-1) & MULT_43(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(17)(MULT_SIZE-1) & MULT_44(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(18)<=signed(MULT_43(18)(MULT_SIZE-1) & MULT_43(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(18)(MULT_SIZE-1) & MULT_44(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(19)<=signed(MULT_43(19)(MULT_SIZE-1) & MULT_43(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(19)(MULT_SIZE-1) & MULT_44(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(20)<=signed(MULT_43(20)(MULT_SIZE-1) & MULT_43(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(20)(MULT_SIZE-1) & MULT_44(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(21)<=signed(MULT_43(21)(MULT_SIZE-1) & MULT_43(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(21)(MULT_SIZE-1) & MULT_44(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(22)<=signed(MULT_43(22)(MULT_SIZE-1) & MULT_43(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(22)(MULT_SIZE-1) & MULT_44(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(23)<=signed(MULT_43(23)(MULT_SIZE-1) & MULT_43(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(23)(MULT_SIZE-1) & MULT_44(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(24)<=signed(MULT_43(24)(MULT_SIZE-1) & MULT_43(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(24)(MULT_SIZE-1) & MULT_44(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(25)<=signed(MULT_43(25)(MULT_SIZE-1) & MULT_43(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(25)(MULT_SIZE-1) & MULT_44(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(26)<=signed(MULT_43(26)(MULT_SIZE-1) & MULT_43(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(26)(MULT_SIZE-1) & MULT_44(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(27)<=signed(MULT_43(27)(MULT_SIZE-1) & MULT_43(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(27)(MULT_SIZE-1) & MULT_44(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(28)<=signed(MULT_43(28)(MULT_SIZE-1) & MULT_43(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(28)(MULT_SIZE-1) & MULT_44(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(29)<=signed(MULT_43(29)(MULT_SIZE-1) & MULT_43(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(29)(MULT_SIZE-1) & MULT_44(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(30)<=signed(MULT_43(30)(MULT_SIZE-1) & MULT_43(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(30)(MULT_SIZE-1) & MULT_44(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(31)<=signed(MULT_43(31)(MULT_SIZE-1) & MULT_43(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(31)(MULT_SIZE-1) & MULT_44(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(32)<=signed(MULT_43(32)(MULT_SIZE-1) & MULT_43(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(32)(MULT_SIZE-1) & MULT_44(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(33)<=signed(MULT_43(33)(MULT_SIZE-1) & MULT_43(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(33)(MULT_SIZE-1) & MULT_44(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(34)<=signed(MULT_43(34)(MULT_SIZE-1) & MULT_43(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(34)(MULT_SIZE-1) & MULT_44(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(35)<=signed(MULT_43(35)(MULT_SIZE-1) & MULT_43(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(35)(MULT_SIZE-1) & MULT_44(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(36)<=signed(MULT_43(36)(MULT_SIZE-1) & MULT_43(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(36)(MULT_SIZE-1) & MULT_44(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(37)<=signed(MULT_43(37)(MULT_SIZE-1) & MULT_43(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(37)(MULT_SIZE-1) & MULT_44(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(38)<=signed(MULT_43(38)(MULT_SIZE-1) & MULT_43(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(38)(MULT_SIZE-1) & MULT_44(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(39)<=signed(MULT_43(39)(MULT_SIZE-1) & MULT_43(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(39)(MULT_SIZE-1) & MULT_44(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(40)<=signed(MULT_43(40)(MULT_SIZE-1) & MULT_43(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(40)(MULT_SIZE-1) & MULT_44(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(41)<=signed(MULT_43(41)(MULT_SIZE-1) & MULT_43(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(41)(MULT_SIZE-1) & MULT_44(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(42)<=signed(MULT_43(42)(MULT_SIZE-1) & MULT_43(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(42)(MULT_SIZE-1) & MULT_44(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(43)<=signed(MULT_43(43)(MULT_SIZE-1) & MULT_43(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(43)(MULT_SIZE-1) & MULT_44(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(44)<=signed(MULT_43(44)(MULT_SIZE-1) & MULT_43(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(44)(MULT_SIZE-1) & MULT_44(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(45)<=signed(MULT_43(45)(MULT_SIZE-1) & MULT_43(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(45)(MULT_SIZE-1) & MULT_44(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(46)<=signed(MULT_43(46)(MULT_SIZE-1) & MULT_43(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(46)(MULT_SIZE-1) & MULT_44(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(47)<=signed(MULT_43(47)(MULT_SIZE-1) & MULT_43(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(47)(MULT_SIZE-1) & MULT_44(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(48)<=signed(MULT_43(48)(MULT_SIZE-1) & MULT_43(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(48)(MULT_SIZE-1) & MULT_44(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(49)<=signed(MULT_43(49)(MULT_SIZE-1) & MULT_43(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(49)(MULT_SIZE-1) & MULT_44(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(50)<=signed(MULT_43(50)(MULT_SIZE-1) & MULT_43(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(50)(MULT_SIZE-1) & MULT_44(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(51)<=signed(MULT_43(51)(MULT_SIZE-1) & MULT_43(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(51)(MULT_SIZE-1) & MULT_44(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(52)<=signed(MULT_43(52)(MULT_SIZE-1) & MULT_43(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(52)(MULT_SIZE-1) & MULT_44(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(53)<=signed(MULT_43(53)(MULT_SIZE-1) & MULT_43(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(53)(MULT_SIZE-1) & MULT_44(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(54)<=signed(MULT_43(54)(MULT_SIZE-1) & MULT_43(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(54)(MULT_SIZE-1) & MULT_44(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(55)<=signed(MULT_43(55)(MULT_SIZE-1) & MULT_43(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(55)(MULT_SIZE-1) & MULT_44(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(56)<=signed(MULT_43(56)(MULT_SIZE-1) & MULT_43(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(56)(MULT_SIZE-1) & MULT_44(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(57)<=signed(MULT_43(57)(MULT_SIZE-1) & MULT_43(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(57)(MULT_SIZE-1) & MULT_44(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(58)<=signed(MULT_43(58)(MULT_SIZE-1) & MULT_43(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(58)(MULT_SIZE-1) & MULT_44(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(59)<=signed(MULT_43(59)(MULT_SIZE-1) & MULT_43(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(59)(MULT_SIZE-1) & MULT_44(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(60)<=signed(MULT_43(60)(MULT_SIZE-1) & MULT_43(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(60)(MULT_SIZE-1) & MULT_44(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(61)<=signed(MULT_43(61)(MULT_SIZE-1) & MULT_43(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(61)(MULT_SIZE-1) & MULT_44(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(62)<=signed(MULT_43(62)(MULT_SIZE-1) & MULT_43(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(62)(MULT_SIZE-1) & MULT_44(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(63)<=signed(MULT_43(63)(MULT_SIZE-1) & MULT_43(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(63)(MULT_SIZE-1) & MULT_44(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(64)<=signed(MULT_43(64)(MULT_SIZE-1) & MULT_43(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(64)(MULT_SIZE-1) & MULT_44(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(65)<=signed(MULT_43(65)(MULT_SIZE-1) & MULT_43(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(65)(MULT_SIZE-1) & MULT_44(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(66)<=signed(MULT_43(66)(MULT_SIZE-1) & MULT_43(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(66)(MULT_SIZE-1) & MULT_44(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(67)<=signed(MULT_43(67)(MULT_SIZE-1) & MULT_43(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(67)(MULT_SIZE-1) & MULT_44(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(68)<=signed(MULT_43(68)(MULT_SIZE-1) & MULT_43(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(68)(MULT_SIZE-1) & MULT_44(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(69)<=signed(MULT_43(69)(MULT_SIZE-1) & MULT_43(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(69)(MULT_SIZE-1) & MULT_44(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(70)<=signed(MULT_43(70)(MULT_SIZE-1) & MULT_43(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(70)(MULT_SIZE-1) & MULT_44(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(71)<=signed(MULT_43(71)(MULT_SIZE-1) & MULT_43(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(71)(MULT_SIZE-1) & MULT_44(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(72)<=signed(MULT_43(72)(MULT_SIZE-1) & MULT_43(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(72)(MULT_SIZE-1) & MULT_44(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(73)<=signed(MULT_43(73)(MULT_SIZE-1) & MULT_43(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(73)(MULT_SIZE-1) & MULT_44(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(74)<=signed(MULT_43(74)(MULT_SIZE-1) & MULT_43(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(74)(MULT_SIZE-1) & MULT_44(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(75)<=signed(MULT_43(75)(MULT_SIZE-1) & MULT_43(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(75)(MULT_SIZE-1) & MULT_44(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(76)<=signed(MULT_43(76)(MULT_SIZE-1) & MULT_43(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(76)(MULT_SIZE-1) & MULT_44(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(77)<=signed(MULT_43(77)(MULT_SIZE-1) & MULT_43(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(77)(MULT_SIZE-1) & MULT_44(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(78)<=signed(MULT_43(78)(MULT_SIZE-1) & MULT_43(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(78)(MULT_SIZE-1) & MULT_44(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(79)<=signed(MULT_43(79)(MULT_SIZE-1) & MULT_43(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(79)(MULT_SIZE-1) & MULT_44(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(80)<=signed(MULT_43(80)(MULT_SIZE-1) & MULT_43(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(80)(MULT_SIZE-1) & MULT_44(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(81)<=signed(MULT_43(81)(MULT_SIZE-1) & MULT_43(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(81)(MULT_SIZE-1) & MULT_44(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(82)<=signed(MULT_43(82)(MULT_SIZE-1) & MULT_43(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(82)(MULT_SIZE-1) & MULT_44(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_22(83)<=signed(MULT_43(83)(MULT_SIZE-1) & MULT_43(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_44(83)(MULT_SIZE-1) & MULT_44(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_23(0)<=signed(MULT_45(0)(MULT_SIZE-1) & MULT_45(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(0)(MULT_SIZE-1) & MULT_46(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(1)<=signed(MULT_45(1)(MULT_SIZE-1) & MULT_45(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(1)(MULT_SIZE-1) & MULT_46(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(2)<=signed(MULT_45(2)(MULT_SIZE-1) & MULT_45(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(2)(MULT_SIZE-1) & MULT_46(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(3)<=signed(MULT_45(3)(MULT_SIZE-1) & MULT_45(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(3)(MULT_SIZE-1) & MULT_46(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(4)<=signed(MULT_45(4)(MULT_SIZE-1) & MULT_45(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(4)(MULT_SIZE-1) & MULT_46(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(5)<=signed(MULT_45(5)(MULT_SIZE-1) & MULT_45(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(5)(MULT_SIZE-1) & MULT_46(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(6)<=signed(MULT_45(6)(MULT_SIZE-1) & MULT_45(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(6)(MULT_SIZE-1) & MULT_46(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(7)<=signed(MULT_45(7)(MULT_SIZE-1) & MULT_45(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(7)(MULT_SIZE-1) & MULT_46(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(8)<=signed(MULT_45(8)(MULT_SIZE-1) & MULT_45(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(8)(MULT_SIZE-1) & MULT_46(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(9)<=signed(MULT_45(9)(MULT_SIZE-1) & MULT_45(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(9)(MULT_SIZE-1) & MULT_46(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(10)<=signed(MULT_45(10)(MULT_SIZE-1) & MULT_45(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(10)(MULT_SIZE-1) & MULT_46(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(11)<=signed(MULT_45(11)(MULT_SIZE-1) & MULT_45(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(11)(MULT_SIZE-1) & MULT_46(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(12)<=signed(MULT_45(12)(MULT_SIZE-1) & MULT_45(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(12)(MULT_SIZE-1) & MULT_46(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(13)<=signed(MULT_45(13)(MULT_SIZE-1) & MULT_45(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(13)(MULT_SIZE-1) & MULT_46(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(14)<=signed(MULT_45(14)(MULT_SIZE-1) & MULT_45(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(14)(MULT_SIZE-1) & MULT_46(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(15)<=signed(MULT_45(15)(MULT_SIZE-1) & MULT_45(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(15)(MULT_SIZE-1) & MULT_46(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(16)<=signed(MULT_45(16)(MULT_SIZE-1) & MULT_45(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(16)(MULT_SIZE-1) & MULT_46(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(17)<=signed(MULT_45(17)(MULT_SIZE-1) & MULT_45(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(17)(MULT_SIZE-1) & MULT_46(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(18)<=signed(MULT_45(18)(MULT_SIZE-1) & MULT_45(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(18)(MULT_SIZE-1) & MULT_46(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(19)<=signed(MULT_45(19)(MULT_SIZE-1) & MULT_45(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(19)(MULT_SIZE-1) & MULT_46(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(20)<=signed(MULT_45(20)(MULT_SIZE-1) & MULT_45(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(20)(MULT_SIZE-1) & MULT_46(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(21)<=signed(MULT_45(21)(MULT_SIZE-1) & MULT_45(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(21)(MULT_SIZE-1) & MULT_46(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(22)<=signed(MULT_45(22)(MULT_SIZE-1) & MULT_45(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(22)(MULT_SIZE-1) & MULT_46(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(23)<=signed(MULT_45(23)(MULT_SIZE-1) & MULT_45(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(23)(MULT_SIZE-1) & MULT_46(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(24)<=signed(MULT_45(24)(MULT_SIZE-1) & MULT_45(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(24)(MULT_SIZE-1) & MULT_46(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(25)<=signed(MULT_45(25)(MULT_SIZE-1) & MULT_45(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(25)(MULT_SIZE-1) & MULT_46(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(26)<=signed(MULT_45(26)(MULT_SIZE-1) & MULT_45(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(26)(MULT_SIZE-1) & MULT_46(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(27)<=signed(MULT_45(27)(MULT_SIZE-1) & MULT_45(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(27)(MULT_SIZE-1) & MULT_46(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(28)<=signed(MULT_45(28)(MULT_SIZE-1) & MULT_45(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(28)(MULT_SIZE-1) & MULT_46(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(29)<=signed(MULT_45(29)(MULT_SIZE-1) & MULT_45(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(29)(MULT_SIZE-1) & MULT_46(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(30)<=signed(MULT_45(30)(MULT_SIZE-1) & MULT_45(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(30)(MULT_SIZE-1) & MULT_46(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(31)<=signed(MULT_45(31)(MULT_SIZE-1) & MULT_45(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(31)(MULT_SIZE-1) & MULT_46(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(32)<=signed(MULT_45(32)(MULT_SIZE-1) & MULT_45(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(32)(MULT_SIZE-1) & MULT_46(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(33)<=signed(MULT_45(33)(MULT_SIZE-1) & MULT_45(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(33)(MULT_SIZE-1) & MULT_46(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(34)<=signed(MULT_45(34)(MULT_SIZE-1) & MULT_45(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(34)(MULT_SIZE-1) & MULT_46(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(35)<=signed(MULT_45(35)(MULT_SIZE-1) & MULT_45(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(35)(MULT_SIZE-1) & MULT_46(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(36)<=signed(MULT_45(36)(MULT_SIZE-1) & MULT_45(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(36)(MULT_SIZE-1) & MULT_46(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(37)<=signed(MULT_45(37)(MULT_SIZE-1) & MULT_45(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(37)(MULT_SIZE-1) & MULT_46(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(38)<=signed(MULT_45(38)(MULT_SIZE-1) & MULT_45(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(38)(MULT_SIZE-1) & MULT_46(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(39)<=signed(MULT_45(39)(MULT_SIZE-1) & MULT_45(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(39)(MULT_SIZE-1) & MULT_46(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(40)<=signed(MULT_45(40)(MULT_SIZE-1) & MULT_45(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(40)(MULT_SIZE-1) & MULT_46(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(41)<=signed(MULT_45(41)(MULT_SIZE-1) & MULT_45(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(41)(MULT_SIZE-1) & MULT_46(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(42)<=signed(MULT_45(42)(MULT_SIZE-1) & MULT_45(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(42)(MULT_SIZE-1) & MULT_46(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(43)<=signed(MULT_45(43)(MULT_SIZE-1) & MULT_45(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(43)(MULT_SIZE-1) & MULT_46(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(44)<=signed(MULT_45(44)(MULT_SIZE-1) & MULT_45(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(44)(MULT_SIZE-1) & MULT_46(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(45)<=signed(MULT_45(45)(MULT_SIZE-1) & MULT_45(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(45)(MULT_SIZE-1) & MULT_46(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(46)<=signed(MULT_45(46)(MULT_SIZE-1) & MULT_45(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(46)(MULT_SIZE-1) & MULT_46(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(47)<=signed(MULT_45(47)(MULT_SIZE-1) & MULT_45(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(47)(MULT_SIZE-1) & MULT_46(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(48)<=signed(MULT_45(48)(MULT_SIZE-1) & MULT_45(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(48)(MULT_SIZE-1) & MULT_46(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(49)<=signed(MULT_45(49)(MULT_SIZE-1) & MULT_45(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(49)(MULT_SIZE-1) & MULT_46(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(50)<=signed(MULT_45(50)(MULT_SIZE-1) & MULT_45(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(50)(MULT_SIZE-1) & MULT_46(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(51)<=signed(MULT_45(51)(MULT_SIZE-1) & MULT_45(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(51)(MULT_SIZE-1) & MULT_46(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(52)<=signed(MULT_45(52)(MULT_SIZE-1) & MULT_45(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(52)(MULT_SIZE-1) & MULT_46(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(53)<=signed(MULT_45(53)(MULT_SIZE-1) & MULT_45(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(53)(MULT_SIZE-1) & MULT_46(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(54)<=signed(MULT_45(54)(MULT_SIZE-1) & MULT_45(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(54)(MULT_SIZE-1) & MULT_46(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(55)<=signed(MULT_45(55)(MULT_SIZE-1) & MULT_45(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(55)(MULT_SIZE-1) & MULT_46(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(56)<=signed(MULT_45(56)(MULT_SIZE-1) & MULT_45(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(56)(MULT_SIZE-1) & MULT_46(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(57)<=signed(MULT_45(57)(MULT_SIZE-1) & MULT_45(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(57)(MULT_SIZE-1) & MULT_46(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(58)<=signed(MULT_45(58)(MULT_SIZE-1) & MULT_45(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(58)(MULT_SIZE-1) & MULT_46(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(59)<=signed(MULT_45(59)(MULT_SIZE-1) & MULT_45(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(59)(MULT_SIZE-1) & MULT_46(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(60)<=signed(MULT_45(60)(MULT_SIZE-1) & MULT_45(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(60)(MULT_SIZE-1) & MULT_46(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(61)<=signed(MULT_45(61)(MULT_SIZE-1) & MULT_45(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(61)(MULT_SIZE-1) & MULT_46(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(62)<=signed(MULT_45(62)(MULT_SIZE-1) & MULT_45(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(62)(MULT_SIZE-1) & MULT_46(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(63)<=signed(MULT_45(63)(MULT_SIZE-1) & MULT_45(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(63)(MULT_SIZE-1) & MULT_46(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(64)<=signed(MULT_45(64)(MULT_SIZE-1) & MULT_45(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(64)(MULT_SIZE-1) & MULT_46(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(65)<=signed(MULT_45(65)(MULT_SIZE-1) & MULT_45(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(65)(MULT_SIZE-1) & MULT_46(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(66)<=signed(MULT_45(66)(MULT_SIZE-1) & MULT_45(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(66)(MULT_SIZE-1) & MULT_46(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(67)<=signed(MULT_45(67)(MULT_SIZE-1) & MULT_45(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(67)(MULT_SIZE-1) & MULT_46(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(68)<=signed(MULT_45(68)(MULT_SIZE-1) & MULT_45(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(68)(MULT_SIZE-1) & MULT_46(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(69)<=signed(MULT_45(69)(MULT_SIZE-1) & MULT_45(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(69)(MULT_SIZE-1) & MULT_46(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(70)<=signed(MULT_45(70)(MULT_SIZE-1) & MULT_45(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(70)(MULT_SIZE-1) & MULT_46(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(71)<=signed(MULT_45(71)(MULT_SIZE-1) & MULT_45(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(71)(MULT_SIZE-1) & MULT_46(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(72)<=signed(MULT_45(72)(MULT_SIZE-1) & MULT_45(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(72)(MULT_SIZE-1) & MULT_46(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(73)<=signed(MULT_45(73)(MULT_SIZE-1) & MULT_45(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(73)(MULT_SIZE-1) & MULT_46(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(74)<=signed(MULT_45(74)(MULT_SIZE-1) & MULT_45(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(74)(MULT_SIZE-1) & MULT_46(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(75)<=signed(MULT_45(75)(MULT_SIZE-1) & MULT_45(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(75)(MULT_SIZE-1) & MULT_46(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(76)<=signed(MULT_45(76)(MULT_SIZE-1) & MULT_45(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(76)(MULT_SIZE-1) & MULT_46(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(77)<=signed(MULT_45(77)(MULT_SIZE-1) & MULT_45(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(77)(MULT_SIZE-1) & MULT_46(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(78)<=signed(MULT_45(78)(MULT_SIZE-1) & MULT_45(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(78)(MULT_SIZE-1) & MULT_46(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(79)<=signed(MULT_45(79)(MULT_SIZE-1) & MULT_45(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(79)(MULT_SIZE-1) & MULT_46(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(80)<=signed(MULT_45(80)(MULT_SIZE-1) & MULT_45(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(80)(MULT_SIZE-1) & MULT_46(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(81)<=signed(MULT_45(81)(MULT_SIZE-1) & MULT_45(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(81)(MULT_SIZE-1) & MULT_46(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(82)<=signed(MULT_45(82)(MULT_SIZE-1) & MULT_45(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(82)(MULT_SIZE-1) & MULT_46(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_23(83)<=signed(MULT_45(83)(MULT_SIZE-1) & MULT_45(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_46(83)(MULT_SIZE-1) & MULT_46(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_24(0)<=signed(MULT_47(0)(MULT_SIZE-1) & MULT_47(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(0)(MULT_SIZE-1) & MULT_48(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(1)<=signed(MULT_47(1)(MULT_SIZE-1) & MULT_47(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(1)(MULT_SIZE-1) & MULT_48(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(2)<=signed(MULT_47(2)(MULT_SIZE-1) & MULT_47(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(2)(MULT_SIZE-1) & MULT_48(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(3)<=signed(MULT_47(3)(MULT_SIZE-1) & MULT_47(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(3)(MULT_SIZE-1) & MULT_48(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(4)<=signed(MULT_47(4)(MULT_SIZE-1) & MULT_47(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(4)(MULT_SIZE-1) & MULT_48(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(5)<=signed(MULT_47(5)(MULT_SIZE-1) & MULT_47(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(5)(MULT_SIZE-1) & MULT_48(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(6)<=signed(MULT_47(6)(MULT_SIZE-1) & MULT_47(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(6)(MULT_SIZE-1) & MULT_48(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(7)<=signed(MULT_47(7)(MULT_SIZE-1) & MULT_47(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(7)(MULT_SIZE-1) & MULT_48(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(8)<=signed(MULT_47(8)(MULT_SIZE-1) & MULT_47(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(8)(MULT_SIZE-1) & MULT_48(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(9)<=signed(MULT_47(9)(MULT_SIZE-1) & MULT_47(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(9)(MULT_SIZE-1) & MULT_48(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(10)<=signed(MULT_47(10)(MULT_SIZE-1) & MULT_47(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(10)(MULT_SIZE-1) & MULT_48(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(11)<=signed(MULT_47(11)(MULT_SIZE-1) & MULT_47(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(11)(MULT_SIZE-1) & MULT_48(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(12)<=signed(MULT_47(12)(MULT_SIZE-1) & MULT_47(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(12)(MULT_SIZE-1) & MULT_48(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(13)<=signed(MULT_47(13)(MULT_SIZE-1) & MULT_47(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(13)(MULT_SIZE-1) & MULT_48(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(14)<=signed(MULT_47(14)(MULT_SIZE-1) & MULT_47(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(14)(MULT_SIZE-1) & MULT_48(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(15)<=signed(MULT_47(15)(MULT_SIZE-1) & MULT_47(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(15)(MULT_SIZE-1) & MULT_48(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(16)<=signed(MULT_47(16)(MULT_SIZE-1) & MULT_47(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(16)(MULT_SIZE-1) & MULT_48(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(17)<=signed(MULT_47(17)(MULT_SIZE-1) & MULT_47(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(17)(MULT_SIZE-1) & MULT_48(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(18)<=signed(MULT_47(18)(MULT_SIZE-1) & MULT_47(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(18)(MULT_SIZE-1) & MULT_48(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(19)<=signed(MULT_47(19)(MULT_SIZE-1) & MULT_47(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(19)(MULT_SIZE-1) & MULT_48(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(20)<=signed(MULT_47(20)(MULT_SIZE-1) & MULT_47(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(20)(MULT_SIZE-1) & MULT_48(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(21)<=signed(MULT_47(21)(MULT_SIZE-1) & MULT_47(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(21)(MULT_SIZE-1) & MULT_48(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(22)<=signed(MULT_47(22)(MULT_SIZE-1) & MULT_47(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(22)(MULT_SIZE-1) & MULT_48(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(23)<=signed(MULT_47(23)(MULT_SIZE-1) & MULT_47(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(23)(MULT_SIZE-1) & MULT_48(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(24)<=signed(MULT_47(24)(MULT_SIZE-1) & MULT_47(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(24)(MULT_SIZE-1) & MULT_48(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(25)<=signed(MULT_47(25)(MULT_SIZE-1) & MULT_47(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(25)(MULT_SIZE-1) & MULT_48(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(26)<=signed(MULT_47(26)(MULT_SIZE-1) & MULT_47(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(26)(MULT_SIZE-1) & MULT_48(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(27)<=signed(MULT_47(27)(MULT_SIZE-1) & MULT_47(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(27)(MULT_SIZE-1) & MULT_48(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(28)<=signed(MULT_47(28)(MULT_SIZE-1) & MULT_47(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(28)(MULT_SIZE-1) & MULT_48(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(29)<=signed(MULT_47(29)(MULT_SIZE-1) & MULT_47(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(29)(MULT_SIZE-1) & MULT_48(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(30)<=signed(MULT_47(30)(MULT_SIZE-1) & MULT_47(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(30)(MULT_SIZE-1) & MULT_48(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(31)<=signed(MULT_47(31)(MULT_SIZE-1) & MULT_47(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(31)(MULT_SIZE-1) & MULT_48(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(32)<=signed(MULT_47(32)(MULT_SIZE-1) & MULT_47(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(32)(MULT_SIZE-1) & MULT_48(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(33)<=signed(MULT_47(33)(MULT_SIZE-1) & MULT_47(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(33)(MULT_SIZE-1) & MULT_48(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(34)<=signed(MULT_47(34)(MULT_SIZE-1) & MULT_47(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(34)(MULT_SIZE-1) & MULT_48(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(35)<=signed(MULT_47(35)(MULT_SIZE-1) & MULT_47(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(35)(MULT_SIZE-1) & MULT_48(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(36)<=signed(MULT_47(36)(MULT_SIZE-1) & MULT_47(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(36)(MULT_SIZE-1) & MULT_48(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(37)<=signed(MULT_47(37)(MULT_SIZE-1) & MULT_47(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(37)(MULT_SIZE-1) & MULT_48(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(38)<=signed(MULT_47(38)(MULT_SIZE-1) & MULT_47(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(38)(MULT_SIZE-1) & MULT_48(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(39)<=signed(MULT_47(39)(MULT_SIZE-1) & MULT_47(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(39)(MULT_SIZE-1) & MULT_48(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(40)<=signed(MULT_47(40)(MULT_SIZE-1) & MULT_47(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(40)(MULT_SIZE-1) & MULT_48(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(41)<=signed(MULT_47(41)(MULT_SIZE-1) & MULT_47(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(41)(MULT_SIZE-1) & MULT_48(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(42)<=signed(MULT_47(42)(MULT_SIZE-1) & MULT_47(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(42)(MULT_SIZE-1) & MULT_48(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(43)<=signed(MULT_47(43)(MULT_SIZE-1) & MULT_47(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(43)(MULT_SIZE-1) & MULT_48(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(44)<=signed(MULT_47(44)(MULT_SIZE-1) & MULT_47(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(44)(MULT_SIZE-1) & MULT_48(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(45)<=signed(MULT_47(45)(MULT_SIZE-1) & MULT_47(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(45)(MULT_SIZE-1) & MULT_48(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(46)<=signed(MULT_47(46)(MULT_SIZE-1) & MULT_47(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(46)(MULT_SIZE-1) & MULT_48(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(47)<=signed(MULT_47(47)(MULT_SIZE-1) & MULT_47(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(47)(MULT_SIZE-1) & MULT_48(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(48)<=signed(MULT_47(48)(MULT_SIZE-1) & MULT_47(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(48)(MULT_SIZE-1) & MULT_48(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(49)<=signed(MULT_47(49)(MULT_SIZE-1) & MULT_47(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(49)(MULT_SIZE-1) & MULT_48(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(50)<=signed(MULT_47(50)(MULT_SIZE-1) & MULT_47(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(50)(MULT_SIZE-1) & MULT_48(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(51)<=signed(MULT_47(51)(MULT_SIZE-1) & MULT_47(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(51)(MULT_SIZE-1) & MULT_48(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(52)<=signed(MULT_47(52)(MULT_SIZE-1) & MULT_47(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(52)(MULT_SIZE-1) & MULT_48(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(53)<=signed(MULT_47(53)(MULT_SIZE-1) & MULT_47(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(53)(MULT_SIZE-1) & MULT_48(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(54)<=signed(MULT_47(54)(MULT_SIZE-1) & MULT_47(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(54)(MULT_SIZE-1) & MULT_48(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(55)<=signed(MULT_47(55)(MULT_SIZE-1) & MULT_47(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(55)(MULT_SIZE-1) & MULT_48(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(56)<=signed(MULT_47(56)(MULT_SIZE-1) & MULT_47(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(56)(MULT_SIZE-1) & MULT_48(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(57)<=signed(MULT_47(57)(MULT_SIZE-1) & MULT_47(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(57)(MULT_SIZE-1) & MULT_48(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(58)<=signed(MULT_47(58)(MULT_SIZE-1) & MULT_47(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(58)(MULT_SIZE-1) & MULT_48(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(59)<=signed(MULT_47(59)(MULT_SIZE-1) & MULT_47(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(59)(MULT_SIZE-1) & MULT_48(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(60)<=signed(MULT_47(60)(MULT_SIZE-1) & MULT_47(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(60)(MULT_SIZE-1) & MULT_48(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(61)<=signed(MULT_47(61)(MULT_SIZE-1) & MULT_47(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(61)(MULT_SIZE-1) & MULT_48(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(62)<=signed(MULT_47(62)(MULT_SIZE-1) & MULT_47(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(62)(MULT_SIZE-1) & MULT_48(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(63)<=signed(MULT_47(63)(MULT_SIZE-1) & MULT_47(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(63)(MULT_SIZE-1) & MULT_48(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(64)<=signed(MULT_47(64)(MULT_SIZE-1) & MULT_47(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(64)(MULT_SIZE-1) & MULT_48(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(65)<=signed(MULT_47(65)(MULT_SIZE-1) & MULT_47(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(65)(MULT_SIZE-1) & MULT_48(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(66)<=signed(MULT_47(66)(MULT_SIZE-1) & MULT_47(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(66)(MULT_SIZE-1) & MULT_48(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(67)<=signed(MULT_47(67)(MULT_SIZE-1) & MULT_47(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(67)(MULT_SIZE-1) & MULT_48(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(68)<=signed(MULT_47(68)(MULT_SIZE-1) & MULT_47(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(68)(MULT_SIZE-1) & MULT_48(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(69)<=signed(MULT_47(69)(MULT_SIZE-1) & MULT_47(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(69)(MULT_SIZE-1) & MULT_48(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(70)<=signed(MULT_47(70)(MULT_SIZE-1) & MULT_47(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(70)(MULT_SIZE-1) & MULT_48(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(71)<=signed(MULT_47(71)(MULT_SIZE-1) & MULT_47(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(71)(MULT_SIZE-1) & MULT_48(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(72)<=signed(MULT_47(72)(MULT_SIZE-1) & MULT_47(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(72)(MULT_SIZE-1) & MULT_48(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(73)<=signed(MULT_47(73)(MULT_SIZE-1) & MULT_47(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(73)(MULT_SIZE-1) & MULT_48(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(74)<=signed(MULT_47(74)(MULT_SIZE-1) & MULT_47(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(74)(MULT_SIZE-1) & MULT_48(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(75)<=signed(MULT_47(75)(MULT_SIZE-1) & MULT_47(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(75)(MULT_SIZE-1) & MULT_48(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(76)<=signed(MULT_47(76)(MULT_SIZE-1) & MULT_47(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(76)(MULT_SIZE-1) & MULT_48(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(77)<=signed(MULT_47(77)(MULT_SIZE-1) & MULT_47(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(77)(MULT_SIZE-1) & MULT_48(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(78)<=signed(MULT_47(78)(MULT_SIZE-1) & MULT_47(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(78)(MULT_SIZE-1) & MULT_48(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(79)<=signed(MULT_47(79)(MULT_SIZE-1) & MULT_47(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(79)(MULT_SIZE-1) & MULT_48(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(80)<=signed(MULT_47(80)(MULT_SIZE-1) & MULT_47(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(80)(MULT_SIZE-1) & MULT_48(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(81)<=signed(MULT_47(81)(MULT_SIZE-1) & MULT_47(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(81)(MULT_SIZE-1) & MULT_48(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(82)<=signed(MULT_47(82)(MULT_SIZE-1) & MULT_47(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(82)(MULT_SIZE-1) & MULT_48(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_24(83)<=signed(MULT_47(83)(MULT_SIZE-1) & MULT_47(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_48(83)(MULT_SIZE-1) & MULT_48(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_25(0)<=signed(MULT_49(0)(MULT_SIZE-1) & MULT_49(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(0)(MULT_SIZE-1) & MULT_50(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(1)<=signed(MULT_49(1)(MULT_SIZE-1) & MULT_49(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(1)(MULT_SIZE-1) & MULT_50(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(2)<=signed(MULT_49(2)(MULT_SIZE-1) & MULT_49(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(2)(MULT_SIZE-1) & MULT_50(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(3)<=signed(MULT_49(3)(MULT_SIZE-1) & MULT_49(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(3)(MULT_SIZE-1) & MULT_50(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(4)<=signed(MULT_49(4)(MULT_SIZE-1) & MULT_49(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(4)(MULT_SIZE-1) & MULT_50(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(5)<=signed(MULT_49(5)(MULT_SIZE-1) & MULT_49(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(5)(MULT_SIZE-1) & MULT_50(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(6)<=signed(MULT_49(6)(MULT_SIZE-1) & MULT_49(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(6)(MULT_SIZE-1) & MULT_50(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(7)<=signed(MULT_49(7)(MULT_SIZE-1) & MULT_49(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(7)(MULT_SIZE-1) & MULT_50(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(8)<=signed(MULT_49(8)(MULT_SIZE-1) & MULT_49(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(8)(MULT_SIZE-1) & MULT_50(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(9)<=signed(MULT_49(9)(MULT_SIZE-1) & MULT_49(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(9)(MULT_SIZE-1) & MULT_50(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(10)<=signed(MULT_49(10)(MULT_SIZE-1) & MULT_49(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(10)(MULT_SIZE-1) & MULT_50(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(11)<=signed(MULT_49(11)(MULT_SIZE-1) & MULT_49(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(11)(MULT_SIZE-1) & MULT_50(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(12)<=signed(MULT_49(12)(MULT_SIZE-1) & MULT_49(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(12)(MULT_SIZE-1) & MULT_50(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(13)<=signed(MULT_49(13)(MULT_SIZE-1) & MULT_49(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(13)(MULT_SIZE-1) & MULT_50(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(14)<=signed(MULT_49(14)(MULT_SIZE-1) & MULT_49(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(14)(MULT_SIZE-1) & MULT_50(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(15)<=signed(MULT_49(15)(MULT_SIZE-1) & MULT_49(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(15)(MULT_SIZE-1) & MULT_50(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(16)<=signed(MULT_49(16)(MULT_SIZE-1) & MULT_49(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(16)(MULT_SIZE-1) & MULT_50(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(17)<=signed(MULT_49(17)(MULT_SIZE-1) & MULT_49(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(17)(MULT_SIZE-1) & MULT_50(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(18)<=signed(MULT_49(18)(MULT_SIZE-1) & MULT_49(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(18)(MULT_SIZE-1) & MULT_50(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(19)<=signed(MULT_49(19)(MULT_SIZE-1) & MULT_49(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(19)(MULT_SIZE-1) & MULT_50(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(20)<=signed(MULT_49(20)(MULT_SIZE-1) & MULT_49(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(20)(MULT_SIZE-1) & MULT_50(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(21)<=signed(MULT_49(21)(MULT_SIZE-1) & MULT_49(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(21)(MULT_SIZE-1) & MULT_50(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(22)<=signed(MULT_49(22)(MULT_SIZE-1) & MULT_49(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(22)(MULT_SIZE-1) & MULT_50(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(23)<=signed(MULT_49(23)(MULT_SIZE-1) & MULT_49(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(23)(MULT_SIZE-1) & MULT_50(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(24)<=signed(MULT_49(24)(MULT_SIZE-1) & MULT_49(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(24)(MULT_SIZE-1) & MULT_50(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(25)<=signed(MULT_49(25)(MULT_SIZE-1) & MULT_49(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(25)(MULT_SIZE-1) & MULT_50(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(26)<=signed(MULT_49(26)(MULT_SIZE-1) & MULT_49(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(26)(MULT_SIZE-1) & MULT_50(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(27)<=signed(MULT_49(27)(MULT_SIZE-1) & MULT_49(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(27)(MULT_SIZE-1) & MULT_50(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(28)<=signed(MULT_49(28)(MULT_SIZE-1) & MULT_49(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(28)(MULT_SIZE-1) & MULT_50(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(29)<=signed(MULT_49(29)(MULT_SIZE-1) & MULT_49(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(29)(MULT_SIZE-1) & MULT_50(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(30)<=signed(MULT_49(30)(MULT_SIZE-1) & MULT_49(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(30)(MULT_SIZE-1) & MULT_50(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(31)<=signed(MULT_49(31)(MULT_SIZE-1) & MULT_49(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(31)(MULT_SIZE-1) & MULT_50(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(32)<=signed(MULT_49(32)(MULT_SIZE-1) & MULT_49(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(32)(MULT_SIZE-1) & MULT_50(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(33)<=signed(MULT_49(33)(MULT_SIZE-1) & MULT_49(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(33)(MULT_SIZE-1) & MULT_50(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(34)<=signed(MULT_49(34)(MULT_SIZE-1) & MULT_49(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(34)(MULT_SIZE-1) & MULT_50(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(35)<=signed(MULT_49(35)(MULT_SIZE-1) & MULT_49(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(35)(MULT_SIZE-1) & MULT_50(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(36)<=signed(MULT_49(36)(MULT_SIZE-1) & MULT_49(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(36)(MULT_SIZE-1) & MULT_50(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(37)<=signed(MULT_49(37)(MULT_SIZE-1) & MULT_49(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(37)(MULT_SIZE-1) & MULT_50(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(38)<=signed(MULT_49(38)(MULT_SIZE-1) & MULT_49(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(38)(MULT_SIZE-1) & MULT_50(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(39)<=signed(MULT_49(39)(MULT_SIZE-1) & MULT_49(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(39)(MULT_SIZE-1) & MULT_50(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(40)<=signed(MULT_49(40)(MULT_SIZE-1) & MULT_49(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(40)(MULT_SIZE-1) & MULT_50(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(41)<=signed(MULT_49(41)(MULT_SIZE-1) & MULT_49(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(41)(MULT_SIZE-1) & MULT_50(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(42)<=signed(MULT_49(42)(MULT_SIZE-1) & MULT_49(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(42)(MULT_SIZE-1) & MULT_50(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(43)<=signed(MULT_49(43)(MULT_SIZE-1) & MULT_49(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(43)(MULT_SIZE-1) & MULT_50(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(44)<=signed(MULT_49(44)(MULT_SIZE-1) & MULT_49(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(44)(MULT_SIZE-1) & MULT_50(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(45)<=signed(MULT_49(45)(MULT_SIZE-1) & MULT_49(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(45)(MULT_SIZE-1) & MULT_50(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(46)<=signed(MULT_49(46)(MULT_SIZE-1) & MULT_49(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(46)(MULT_SIZE-1) & MULT_50(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(47)<=signed(MULT_49(47)(MULT_SIZE-1) & MULT_49(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(47)(MULT_SIZE-1) & MULT_50(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(48)<=signed(MULT_49(48)(MULT_SIZE-1) & MULT_49(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(48)(MULT_SIZE-1) & MULT_50(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(49)<=signed(MULT_49(49)(MULT_SIZE-1) & MULT_49(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(49)(MULT_SIZE-1) & MULT_50(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(50)<=signed(MULT_49(50)(MULT_SIZE-1) & MULT_49(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(50)(MULT_SIZE-1) & MULT_50(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(51)<=signed(MULT_49(51)(MULT_SIZE-1) & MULT_49(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(51)(MULT_SIZE-1) & MULT_50(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(52)<=signed(MULT_49(52)(MULT_SIZE-1) & MULT_49(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(52)(MULT_SIZE-1) & MULT_50(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(53)<=signed(MULT_49(53)(MULT_SIZE-1) & MULT_49(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(53)(MULT_SIZE-1) & MULT_50(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(54)<=signed(MULT_49(54)(MULT_SIZE-1) & MULT_49(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(54)(MULT_SIZE-1) & MULT_50(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(55)<=signed(MULT_49(55)(MULT_SIZE-1) & MULT_49(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(55)(MULT_SIZE-1) & MULT_50(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(56)<=signed(MULT_49(56)(MULT_SIZE-1) & MULT_49(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(56)(MULT_SIZE-1) & MULT_50(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(57)<=signed(MULT_49(57)(MULT_SIZE-1) & MULT_49(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(57)(MULT_SIZE-1) & MULT_50(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(58)<=signed(MULT_49(58)(MULT_SIZE-1) & MULT_49(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(58)(MULT_SIZE-1) & MULT_50(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(59)<=signed(MULT_49(59)(MULT_SIZE-1) & MULT_49(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(59)(MULT_SIZE-1) & MULT_50(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(60)<=signed(MULT_49(60)(MULT_SIZE-1) & MULT_49(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(60)(MULT_SIZE-1) & MULT_50(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(61)<=signed(MULT_49(61)(MULT_SIZE-1) & MULT_49(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(61)(MULT_SIZE-1) & MULT_50(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(62)<=signed(MULT_49(62)(MULT_SIZE-1) & MULT_49(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(62)(MULT_SIZE-1) & MULT_50(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(63)<=signed(MULT_49(63)(MULT_SIZE-1) & MULT_49(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(63)(MULT_SIZE-1) & MULT_50(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(64)<=signed(MULT_49(64)(MULT_SIZE-1) & MULT_49(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(64)(MULT_SIZE-1) & MULT_50(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(65)<=signed(MULT_49(65)(MULT_SIZE-1) & MULT_49(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(65)(MULT_SIZE-1) & MULT_50(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(66)<=signed(MULT_49(66)(MULT_SIZE-1) & MULT_49(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(66)(MULT_SIZE-1) & MULT_50(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(67)<=signed(MULT_49(67)(MULT_SIZE-1) & MULT_49(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(67)(MULT_SIZE-1) & MULT_50(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(68)<=signed(MULT_49(68)(MULT_SIZE-1) & MULT_49(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(68)(MULT_SIZE-1) & MULT_50(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(69)<=signed(MULT_49(69)(MULT_SIZE-1) & MULT_49(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(69)(MULT_SIZE-1) & MULT_50(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(70)<=signed(MULT_49(70)(MULT_SIZE-1) & MULT_49(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(70)(MULT_SIZE-1) & MULT_50(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(71)<=signed(MULT_49(71)(MULT_SIZE-1) & MULT_49(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(71)(MULT_SIZE-1) & MULT_50(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(72)<=signed(MULT_49(72)(MULT_SIZE-1) & MULT_49(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(72)(MULT_SIZE-1) & MULT_50(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(73)<=signed(MULT_49(73)(MULT_SIZE-1) & MULT_49(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(73)(MULT_SIZE-1) & MULT_50(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(74)<=signed(MULT_49(74)(MULT_SIZE-1) & MULT_49(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(74)(MULT_SIZE-1) & MULT_50(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(75)<=signed(MULT_49(75)(MULT_SIZE-1) & MULT_49(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(75)(MULT_SIZE-1) & MULT_50(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(76)<=signed(MULT_49(76)(MULT_SIZE-1) & MULT_49(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(76)(MULT_SIZE-1) & MULT_50(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(77)<=signed(MULT_49(77)(MULT_SIZE-1) & MULT_49(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(77)(MULT_SIZE-1) & MULT_50(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(78)<=signed(MULT_49(78)(MULT_SIZE-1) & MULT_49(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(78)(MULT_SIZE-1) & MULT_50(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(79)<=signed(MULT_49(79)(MULT_SIZE-1) & MULT_49(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(79)(MULT_SIZE-1) & MULT_50(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(80)<=signed(MULT_49(80)(MULT_SIZE-1) & MULT_49(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(80)(MULT_SIZE-1) & MULT_50(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(81)<=signed(MULT_49(81)(MULT_SIZE-1) & MULT_49(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(81)(MULT_SIZE-1) & MULT_50(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(82)<=signed(MULT_49(82)(MULT_SIZE-1) & MULT_49(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(82)(MULT_SIZE-1) & MULT_50(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_25(83)<=signed(MULT_49(83)(MULT_SIZE-1) & MULT_49(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_50(83)(MULT_SIZE-1) & MULT_50(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_26(0)<=signed(MULT_51(0)(MULT_SIZE-1) & MULT_51(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(0)(MULT_SIZE-1) & MULT_52(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(1)<=signed(MULT_51(1)(MULT_SIZE-1) & MULT_51(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(1)(MULT_SIZE-1) & MULT_52(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(2)<=signed(MULT_51(2)(MULT_SIZE-1) & MULT_51(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(2)(MULT_SIZE-1) & MULT_52(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(3)<=signed(MULT_51(3)(MULT_SIZE-1) & MULT_51(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(3)(MULT_SIZE-1) & MULT_52(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(4)<=signed(MULT_51(4)(MULT_SIZE-1) & MULT_51(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(4)(MULT_SIZE-1) & MULT_52(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(5)<=signed(MULT_51(5)(MULT_SIZE-1) & MULT_51(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(5)(MULT_SIZE-1) & MULT_52(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(6)<=signed(MULT_51(6)(MULT_SIZE-1) & MULT_51(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(6)(MULT_SIZE-1) & MULT_52(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(7)<=signed(MULT_51(7)(MULT_SIZE-1) & MULT_51(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(7)(MULT_SIZE-1) & MULT_52(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(8)<=signed(MULT_51(8)(MULT_SIZE-1) & MULT_51(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(8)(MULT_SIZE-1) & MULT_52(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(9)<=signed(MULT_51(9)(MULT_SIZE-1) & MULT_51(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(9)(MULT_SIZE-1) & MULT_52(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(10)<=signed(MULT_51(10)(MULT_SIZE-1) & MULT_51(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(10)(MULT_SIZE-1) & MULT_52(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(11)<=signed(MULT_51(11)(MULT_SIZE-1) & MULT_51(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(11)(MULT_SIZE-1) & MULT_52(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(12)<=signed(MULT_51(12)(MULT_SIZE-1) & MULT_51(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(12)(MULT_SIZE-1) & MULT_52(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(13)<=signed(MULT_51(13)(MULT_SIZE-1) & MULT_51(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(13)(MULT_SIZE-1) & MULT_52(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(14)<=signed(MULT_51(14)(MULT_SIZE-1) & MULT_51(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(14)(MULT_SIZE-1) & MULT_52(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(15)<=signed(MULT_51(15)(MULT_SIZE-1) & MULT_51(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(15)(MULT_SIZE-1) & MULT_52(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(16)<=signed(MULT_51(16)(MULT_SIZE-1) & MULT_51(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(16)(MULT_SIZE-1) & MULT_52(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(17)<=signed(MULT_51(17)(MULT_SIZE-1) & MULT_51(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(17)(MULT_SIZE-1) & MULT_52(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(18)<=signed(MULT_51(18)(MULT_SIZE-1) & MULT_51(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(18)(MULT_SIZE-1) & MULT_52(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(19)<=signed(MULT_51(19)(MULT_SIZE-1) & MULT_51(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(19)(MULT_SIZE-1) & MULT_52(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(20)<=signed(MULT_51(20)(MULT_SIZE-1) & MULT_51(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(20)(MULT_SIZE-1) & MULT_52(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(21)<=signed(MULT_51(21)(MULT_SIZE-1) & MULT_51(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(21)(MULT_SIZE-1) & MULT_52(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(22)<=signed(MULT_51(22)(MULT_SIZE-1) & MULT_51(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(22)(MULT_SIZE-1) & MULT_52(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(23)<=signed(MULT_51(23)(MULT_SIZE-1) & MULT_51(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(23)(MULT_SIZE-1) & MULT_52(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(24)<=signed(MULT_51(24)(MULT_SIZE-1) & MULT_51(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(24)(MULT_SIZE-1) & MULT_52(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(25)<=signed(MULT_51(25)(MULT_SIZE-1) & MULT_51(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(25)(MULT_SIZE-1) & MULT_52(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(26)<=signed(MULT_51(26)(MULT_SIZE-1) & MULT_51(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(26)(MULT_SIZE-1) & MULT_52(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(27)<=signed(MULT_51(27)(MULT_SIZE-1) & MULT_51(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(27)(MULT_SIZE-1) & MULT_52(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(28)<=signed(MULT_51(28)(MULT_SIZE-1) & MULT_51(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(28)(MULT_SIZE-1) & MULT_52(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(29)<=signed(MULT_51(29)(MULT_SIZE-1) & MULT_51(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(29)(MULT_SIZE-1) & MULT_52(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(30)<=signed(MULT_51(30)(MULT_SIZE-1) & MULT_51(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(30)(MULT_SIZE-1) & MULT_52(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(31)<=signed(MULT_51(31)(MULT_SIZE-1) & MULT_51(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(31)(MULT_SIZE-1) & MULT_52(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(32)<=signed(MULT_51(32)(MULT_SIZE-1) & MULT_51(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(32)(MULT_SIZE-1) & MULT_52(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(33)<=signed(MULT_51(33)(MULT_SIZE-1) & MULT_51(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(33)(MULT_SIZE-1) & MULT_52(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(34)<=signed(MULT_51(34)(MULT_SIZE-1) & MULT_51(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(34)(MULT_SIZE-1) & MULT_52(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(35)<=signed(MULT_51(35)(MULT_SIZE-1) & MULT_51(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(35)(MULT_SIZE-1) & MULT_52(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(36)<=signed(MULT_51(36)(MULT_SIZE-1) & MULT_51(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(36)(MULT_SIZE-1) & MULT_52(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(37)<=signed(MULT_51(37)(MULT_SIZE-1) & MULT_51(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(37)(MULT_SIZE-1) & MULT_52(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(38)<=signed(MULT_51(38)(MULT_SIZE-1) & MULT_51(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(38)(MULT_SIZE-1) & MULT_52(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(39)<=signed(MULT_51(39)(MULT_SIZE-1) & MULT_51(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(39)(MULT_SIZE-1) & MULT_52(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(40)<=signed(MULT_51(40)(MULT_SIZE-1) & MULT_51(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(40)(MULT_SIZE-1) & MULT_52(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(41)<=signed(MULT_51(41)(MULT_SIZE-1) & MULT_51(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(41)(MULT_SIZE-1) & MULT_52(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(42)<=signed(MULT_51(42)(MULT_SIZE-1) & MULT_51(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(42)(MULT_SIZE-1) & MULT_52(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(43)<=signed(MULT_51(43)(MULT_SIZE-1) & MULT_51(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(43)(MULT_SIZE-1) & MULT_52(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(44)<=signed(MULT_51(44)(MULT_SIZE-1) & MULT_51(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(44)(MULT_SIZE-1) & MULT_52(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(45)<=signed(MULT_51(45)(MULT_SIZE-1) & MULT_51(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(45)(MULT_SIZE-1) & MULT_52(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(46)<=signed(MULT_51(46)(MULT_SIZE-1) & MULT_51(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(46)(MULT_SIZE-1) & MULT_52(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(47)<=signed(MULT_51(47)(MULT_SIZE-1) & MULT_51(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(47)(MULT_SIZE-1) & MULT_52(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(48)<=signed(MULT_51(48)(MULT_SIZE-1) & MULT_51(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(48)(MULT_SIZE-1) & MULT_52(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(49)<=signed(MULT_51(49)(MULT_SIZE-1) & MULT_51(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(49)(MULT_SIZE-1) & MULT_52(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(50)<=signed(MULT_51(50)(MULT_SIZE-1) & MULT_51(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(50)(MULT_SIZE-1) & MULT_52(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(51)<=signed(MULT_51(51)(MULT_SIZE-1) & MULT_51(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(51)(MULT_SIZE-1) & MULT_52(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(52)<=signed(MULT_51(52)(MULT_SIZE-1) & MULT_51(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(52)(MULT_SIZE-1) & MULT_52(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(53)<=signed(MULT_51(53)(MULT_SIZE-1) & MULT_51(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(53)(MULT_SIZE-1) & MULT_52(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(54)<=signed(MULT_51(54)(MULT_SIZE-1) & MULT_51(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(54)(MULT_SIZE-1) & MULT_52(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(55)<=signed(MULT_51(55)(MULT_SIZE-1) & MULT_51(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(55)(MULT_SIZE-1) & MULT_52(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(56)<=signed(MULT_51(56)(MULT_SIZE-1) & MULT_51(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(56)(MULT_SIZE-1) & MULT_52(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(57)<=signed(MULT_51(57)(MULT_SIZE-1) & MULT_51(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(57)(MULT_SIZE-1) & MULT_52(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(58)<=signed(MULT_51(58)(MULT_SIZE-1) & MULT_51(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(58)(MULT_SIZE-1) & MULT_52(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(59)<=signed(MULT_51(59)(MULT_SIZE-1) & MULT_51(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(59)(MULT_SIZE-1) & MULT_52(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(60)<=signed(MULT_51(60)(MULT_SIZE-1) & MULT_51(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(60)(MULT_SIZE-1) & MULT_52(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(61)<=signed(MULT_51(61)(MULT_SIZE-1) & MULT_51(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(61)(MULT_SIZE-1) & MULT_52(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(62)<=signed(MULT_51(62)(MULT_SIZE-1) & MULT_51(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(62)(MULT_SIZE-1) & MULT_52(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(63)<=signed(MULT_51(63)(MULT_SIZE-1) & MULT_51(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(63)(MULT_SIZE-1) & MULT_52(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(64)<=signed(MULT_51(64)(MULT_SIZE-1) & MULT_51(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(64)(MULT_SIZE-1) & MULT_52(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(65)<=signed(MULT_51(65)(MULT_SIZE-1) & MULT_51(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(65)(MULT_SIZE-1) & MULT_52(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(66)<=signed(MULT_51(66)(MULT_SIZE-1) & MULT_51(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(66)(MULT_SIZE-1) & MULT_52(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(67)<=signed(MULT_51(67)(MULT_SIZE-1) & MULT_51(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(67)(MULT_SIZE-1) & MULT_52(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(68)<=signed(MULT_51(68)(MULT_SIZE-1) & MULT_51(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(68)(MULT_SIZE-1) & MULT_52(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(69)<=signed(MULT_51(69)(MULT_SIZE-1) & MULT_51(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(69)(MULT_SIZE-1) & MULT_52(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(70)<=signed(MULT_51(70)(MULT_SIZE-1) & MULT_51(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(70)(MULT_SIZE-1) & MULT_52(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(71)<=signed(MULT_51(71)(MULT_SIZE-1) & MULT_51(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(71)(MULT_SIZE-1) & MULT_52(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(72)<=signed(MULT_51(72)(MULT_SIZE-1) & MULT_51(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(72)(MULT_SIZE-1) & MULT_52(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(73)<=signed(MULT_51(73)(MULT_SIZE-1) & MULT_51(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(73)(MULT_SIZE-1) & MULT_52(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(74)<=signed(MULT_51(74)(MULT_SIZE-1) & MULT_51(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(74)(MULT_SIZE-1) & MULT_52(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(75)<=signed(MULT_51(75)(MULT_SIZE-1) & MULT_51(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(75)(MULT_SIZE-1) & MULT_52(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(76)<=signed(MULT_51(76)(MULT_SIZE-1) & MULT_51(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(76)(MULT_SIZE-1) & MULT_52(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(77)<=signed(MULT_51(77)(MULT_SIZE-1) & MULT_51(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(77)(MULT_SIZE-1) & MULT_52(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(78)<=signed(MULT_51(78)(MULT_SIZE-1) & MULT_51(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(78)(MULT_SIZE-1) & MULT_52(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(79)<=signed(MULT_51(79)(MULT_SIZE-1) & MULT_51(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(79)(MULT_SIZE-1) & MULT_52(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(80)<=signed(MULT_51(80)(MULT_SIZE-1) & MULT_51(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(80)(MULT_SIZE-1) & MULT_52(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(81)<=signed(MULT_51(81)(MULT_SIZE-1) & MULT_51(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(81)(MULT_SIZE-1) & MULT_52(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(82)<=signed(MULT_51(82)(MULT_SIZE-1) & MULT_51(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(82)(MULT_SIZE-1) & MULT_52(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_26(83)<=signed(MULT_51(83)(MULT_SIZE-1) & MULT_51(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_52(83)(MULT_SIZE-1) & MULT_52(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_27(0)<=signed(MULT_53(0)(MULT_SIZE-1) & MULT_53(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(0)(MULT_SIZE-1) & MULT_54(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(1)<=signed(MULT_53(1)(MULT_SIZE-1) & MULT_53(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(1)(MULT_SIZE-1) & MULT_54(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(2)<=signed(MULT_53(2)(MULT_SIZE-1) & MULT_53(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(2)(MULT_SIZE-1) & MULT_54(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(3)<=signed(MULT_53(3)(MULT_SIZE-1) & MULT_53(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(3)(MULT_SIZE-1) & MULT_54(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(4)<=signed(MULT_53(4)(MULT_SIZE-1) & MULT_53(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(4)(MULT_SIZE-1) & MULT_54(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(5)<=signed(MULT_53(5)(MULT_SIZE-1) & MULT_53(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(5)(MULT_SIZE-1) & MULT_54(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(6)<=signed(MULT_53(6)(MULT_SIZE-1) & MULT_53(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(6)(MULT_SIZE-1) & MULT_54(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(7)<=signed(MULT_53(7)(MULT_SIZE-1) & MULT_53(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(7)(MULT_SIZE-1) & MULT_54(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(8)<=signed(MULT_53(8)(MULT_SIZE-1) & MULT_53(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(8)(MULT_SIZE-1) & MULT_54(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(9)<=signed(MULT_53(9)(MULT_SIZE-1) & MULT_53(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(9)(MULT_SIZE-1) & MULT_54(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(10)<=signed(MULT_53(10)(MULT_SIZE-1) & MULT_53(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(10)(MULT_SIZE-1) & MULT_54(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(11)<=signed(MULT_53(11)(MULT_SIZE-1) & MULT_53(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(11)(MULT_SIZE-1) & MULT_54(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(12)<=signed(MULT_53(12)(MULT_SIZE-1) & MULT_53(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(12)(MULT_SIZE-1) & MULT_54(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(13)<=signed(MULT_53(13)(MULT_SIZE-1) & MULT_53(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(13)(MULT_SIZE-1) & MULT_54(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(14)<=signed(MULT_53(14)(MULT_SIZE-1) & MULT_53(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(14)(MULT_SIZE-1) & MULT_54(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(15)<=signed(MULT_53(15)(MULT_SIZE-1) & MULT_53(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(15)(MULT_SIZE-1) & MULT_54(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(16)<=signed(MULT_53(16)(MULT_SIZE-1) & MULT_53(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(16)(MULT_SIZE-1) & MULT_54(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(17)<=signed(MULT_53(17)(MULT_SIZE-1) & MULT_53(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(17)(MULT_SIZE-1) & MULT_54(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(18)<=signed(MULT_53(18)(MULT_SIZE-1) & MULT_53(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(18)(MULT_SIZE-1) & MULT_54(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(19)<=signed(MULT_53(19)(MULT_SIZE-1) & MULT_53(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(19)(MULT_SIZE-1) & MULT_54(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(20)<=signed(MULT_53(20)(MULT_SIZE-1) & MULT_53(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(20)(MULT_SIZE-1) & MULT_54(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(21)<=signed(MULT_53(21)(MULT_SIZE-1) & MULT_53(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(21)(MULT_SIZE-1) & MULT_54(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(22)<=signed(MULT_53(22)(MULT_SIZE-1) & MULT_53(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(22)(MULT_SIZE-1) & MULT_54(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(23)<=signed(MULT_53(23)(MULT_SIZE-1) & MULT_53(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(23)(MULT_SIZE-1) & MULT_54(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(24)<=signed(MULT_53(24)(MULT_SIZE-1) & MULT_53(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(24)(MULT_SIZE-1) & MULT_54(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(25)<=signed(MULT_53(25)(MULT_SIZE-1) & MULT_53(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(25)(MULT_SIZE-1) & MULT_54(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(26)<=signed(MULT_53(26)(MULT_SIZE-1) & MULT_53(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(26)(MULT_SIZE-1) & MULT_54(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(27)<=signed(MULT_53(27)(MULT_SIZE-1) & MULT_53(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(27)(MULT_SIZE-1) & MULT_54(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(28)<=signed(MULT_53(28)(MULT_SIZE-1) & MULT_53(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(28)(MULT_SIZE-1) & MULT_54(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(29)<=signed(MULT_53(29)(MULT_SIZE-1) & MULT_53(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(29)(MULT_SIZE-1) & MULT_54(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(30)<=signed(MULT_53(30)(MULT_SIZE-1) & MULT_53(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(30)(MULT_SIZE-1) & MULT_54(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(31)<=signed(MULT_53(31)(MULT_SIZE-1) & MULT_53(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(31)(MULT_SIZE-1) & MULT_54(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(32)<=signed(MULT_53(32)(MULT_SIZE-1) & MULT_53(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(32)(MULT_SIZE-1) & MULT_54(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(33)<=signed(MULT_53(33)(MULT_SIZE-1) & MULT_53(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(33)(MULT_SIZE-1) & MULT_54(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(34)<=signed(MULT_53(34)(MULT_SIZE-1) & MULT_53(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(34)(MULT_SIZE-1) & MULT_54(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(35)<=signed(MULT_53(35)(MULT_SIZE-1) & MULT_53(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(35)(MULT_SIZE-1) & MULT_54(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(36)<=signed(MULT_53(36)(MULT_SIZE-1) & MULT_53(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(36)(MULT_SIZE-1) & MULT_54(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(37)<=signed(MULT_53(37)(MULT_SIZE-1) & MULT_53(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(37)(MULT_SIZE-1) & MULT_54(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(38)<=signed(MULT_53(38)(MULT_SIZE-1) & MULT_53(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(38)(MULT_SIZE-1) & MULT_54(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(39)<=signed(MULT_53(39)(MULT_SIZE-1) & MULT_53(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(39)(MULT_SIZE-1) & MULT_54(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(40)<=signed(MULT_53(40)(MULT_SIZE-1) & MULT_53(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(40)(MULT_SIZE-1) & MULT_54(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(41)<=signed(MULT_53(41)(MULT_SIZE-1) & MULT_53(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(41)(MULT_SIZE-1) & MULT_54(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(42)<=signed(MULT_53(42)(MULT_SIZE-1) & MULT_53(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(42)(MULT_SIZE-1) & MULT_54(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(43)<=signed(MULT_53(43)(MULT_SIZE-1) & MULT_53(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(43)(MULT_SIZE-1) & MULT_54(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(44)<=signed(MULT_53(44)(MULT_SIZE-1) & MULT_53(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(44)(MULT_SIZE-1) & MULT_54(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(45)<=signed(MULT_53(45)(MULT_SIZE-1) & MULT_53(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(45)(MULT_SIZE-1) & MULT_54(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(46)<=signed(MULT_53(46)(MULT_SIZE-1) & MULT_53(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(46)(MULT_SIZE-1) & MULT_54(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(47)<=signed(MULT_53(47)(MULT_SIZE-1) & MULT_53(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(47)(MULT_SIZE-1) & MULT_54(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(48)<=signed(MULT_53(48)(MULT_SIZE-1) & MULT_53(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(48)(MULT_SIZE-1) & MULT_54(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(49)<=signed(MULT_53(49)(MULT_SIZE-1) & MULT_53(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(49)(MULT_SIZE-1) & MULT_54(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(50)<=signed(MULT_53(50)(MULT_SIZE-1) & MULT_53(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(50)(MULT_SIZE-1) & MULT_54(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(51)<=signed(MULT_53(51)(MULT_SIZE-1) & MULT_53(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(51)(MULT_SIZE-1) & MULT_54(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(52)<=signed(MULT_53(52)(MULT_SIZE-1) & MULT_53(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(52)(MULT_SIZE-1) & MULT_54(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(53)<=signed(MULT_53(53)(MULT_SIZE-1) & MULT_53(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(53)(MULT_SIZE-1) & MULT_54(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(54)<=signed(MULT_53(54)(MULT_SIZE-1) & MULT_53(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(54)(MULT_SIZE-1) & MULT_54(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(55)<=signed(MULT_53(55)(MULT_SIZE-1) & MULT_53(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(55)(MULT_SIZE-1) & MULT_54(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(56)<=signed(MULT_53(56)(MULT_SIZE-1) & MULT_53(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(56)(MULT_SIZE-1) & MULT_54(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(57)<=signed(MULT_53(57)(MULT_SIZE-1) & MULT_53(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(57)(MULT_SIZE-1) & MULT_54(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(58)<=signed(MULT_53(58)(MULT_SIZE-1) & MULT_53(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(58)(MULT_SIZE-1) & MULT_54(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(59)<=signed(MULT_53(59)(MULT_SIZE-1) & MULT_53(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(59)(MULT_SIZE-1) & MULT_54(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(60)<=signed(MULT_53(60)(MULT_SIZE-1) & MULT_53(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(60)(MULT_SIZE-1) & MULT_54(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(61)<=signed(MULT_53(61)(MULT_SIZE-1) & MULT_53(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(61)(MULT_SIZE-1) & MULT_54(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(62)<=signed(MULT_53(62)(MULT_SIZE-1) & MULT_53(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(62)(MULT_SIZE-1) & MULT_54(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(63)<=signed(MULT_53(63)(MULT_SIZE-1) & MULT_53(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(63)(MULT_SIZE-1) & MULT_54(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(64)<=signed(MULT_53(64)(MULT_SIZE-1) & MULT_53(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(64)(MULT_SIZE-1) & MULT_54(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(65)<=signed(MULT_53(65)(MULT_SIZE-1) & MULT_53(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(65)(MULT_SIZE-1) & MULT_54(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(66)<=signed(MULT_53(66)(MULT_SIZE-1) & MULT_53(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(66)(MULT_SIZE-1) & MULT_54(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(67)<=signed(MULT_53(67)(MULT_SIZE-1) & MULT_53(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(67)(MULT_SIZE-1) & MULT_54(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(68)<=signed(MULT_53(68)(MULT_SIZE-1) & MULT_53(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(68)(MULT_SIZE-1) & MULT_54(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(69)<=signed(MULT_53(69)(MULT_SIZE-1) & MULT_53(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(69)(MULT_SIZE-1) & MULT_54(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(70)<=signed(MULT_53(70)(MULT_SIZE-1) & MULT_53(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(70)(MULT_SIZE-1) & MULT_54(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(71)<=signed(MULT_53(71)(MULT_SIZE-1) & MULT_53(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(71)(MULT_SIZE-1) & MULT_54(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(72)<=signed(MULT_53(72)(MULT_SIZE-1) & MULT_53(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(72)(MULT_SIZE-1) & MULT_54(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(73)<=signed(MULT_53(73)(MULT_SIZE-1) & MULT_53(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(73)(MULT_SIZE-1) & MULT_54(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(74)<=signed(MULT_53(74)(MULT_SIZE-1) & MULT_53(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(74)(MULT_SIZE-1) & MULT_54(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(75)<=signed(MULT_53(75)(MULT_SIZE-1) & MULT_53(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(75)(MULT_SIZE-1) & MULT_54(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(76)<=signed(MULT_53(76)(MULT_SIZE-1) & MULT_53(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(76)(MULT_SIZE-1) & MULT_54(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(77)<=signed(MULT_53(77)(MULT_SIZE-1) & MULT_53(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(77)(MULT_SIZE-1) & MULT_54(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(78)<=signed(MULT_53(78)(MULT_SIZE-1) & MULT_53(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(78)(MULT_SIZE-1) & MULT_54(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(79)<=signed(MULT_53(79)(MULT_SIZE-1) & MULT_53(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(79)(MULT_SIZE-1) & MULT_54(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(80)<=signed(MULT_53(80)(MULT_SIZE-1) & MULT_53(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(80)(MULT_SIZE-1) & MULT_54(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(81)<=signed(MULT_53(81)(MULT_SIZE-1) & MULT_53(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(81)(MULT_SIZE-1) & MULT_54(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(82)<=signed(MULT_53(82)(MULT_SIZE-1) & MULT_53(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(82)(MULT_SIZE-1) & MULT_54(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_27(83)<=signed(MULT_53(83)(MULT_SIZE-1) & MULT_53(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_54(83)(MULT_SIZE-1) & MULT_54(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_28(0)<=signed(MULT_55(0)(MULT_SIZE-1) & MULT_55(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(0)(MULT_SIZE-1) & MULT_56(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(1)<=signed(MULT_55(1)(MULT_SIZE-1) & MULT_55(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(1)(MULT_SIZE-1) & MULT_56(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(2)<=signed(MULT_55(2)(MULT_SIZE-1) & MULT_55(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(2)(MULT_SIZE-1) & MULT_56(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(3)<=signed(MULT_55(3)(MULT_SIZE-1) & MULT_55(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(3)(MULT_SIZE-1) & MULT_56(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(4)<=signed(MULT_55(4)(MULT_SIZE-1) & MULT_55(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(4)(MULT_SIZE-1) & MULT_56(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(5)<=signed(MULT_55(5)(MULT_SIZE-1) & MULT_55(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(5)(MULT_SIZE-1) & MULT_56(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(6)<=signed(MULT_55(6)(MULT_SIZE-1) & MULT_55(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(6)(MULT_SIZE-1) & MULT_56(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(7)<=signed(MULT_55(7)(MULT_SIZE-1) & MULT_55(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(7)(MULT_SIZE-1) & MULT_56(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(8)<=signed(MULT_55(8)(MULT_SIZE-1) & MULT_55(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(8)(MULT_SIZE-1) & MULT_56(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(9)<=signed(MULT_55(9)(MULT_SIZE-1) & MULT_55(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(9)(MULT_SIZE-1) & MULT_56(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(10)<=signed(MULT_55(10)(MULT_SIZE-1) & MULT_55(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(10)(MULT_SIZE-1) & MULT_56(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(11)<=signed(MULT_55(11)(MULT_SIZE-1) & MULT_55(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(11)(MULT_SIZE-1) & MULT_56(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(12)<=signed(MULT_55(12)(MULT_SIZE-1) & MULT_55(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(12)(MULT_SIZE-1) & MULT_56(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(13)<=signed(MULT_55(13)(MULT_SIZE-1) & MULT_55(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(13)(MULT_SIZE-1) & MULT_56(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(14)<=signed(MULT_55(14)(MULT_SIZE-1) & MULT_55(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(14)(MULT_SIZE-1) & MULT_56(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(15)<=signed(MULT_55(15)(MULT_SIZE-1) & MULT_55(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(15)(MULT_SIZE-1) & MULT_56(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(16)<=signed(MULT_55(16)(MULT_SIZE-1) & MULT_55(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(16)(MULT_SIZE-1) & MULT_56(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(17)<=signed(MULT_55(17)(MULT_SIZE-1) & MULT_55(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(17)(MULT_SIZE-1) & MULT_56(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(18)<=signed(MULT_55(18)(MULT_SIZE-1) & MULT_55(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(18)(MULT_SIZE-1) & MULT_56(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(19)<=signed(MULT_55(19)(MULT_SIZE-1) & MULT_55(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(19)(MULT_SIZE-1) & MULT_56(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(20)<=signed(MULT_55(20)(MULT_SIZE-1) & MULT_55(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(20)(MULT_SIZE-1) & MULT_56(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(21)<=signed(MULT_55(21)(MULT_SIZE-1) & MULT_55(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(21)(MULT_SIZE-1) & MULT_56(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(22)<=signed(MULT_55(22)(MULT_SIZE-1) & MULT_55(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(22)(MULT_SIZE-1) & MULT_56(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(23)<=signed(MULT_55(23)(MULT_SIZE-1) & MULT_55(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(23)(MULT_SIZE-1) & MULT_56(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(24)<=signed(MULT_55(24)(MULT_SIZE-1) & MULT_55(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(24)(MULT_SIZE-1) & MULT_56(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(25)<=signed(MULT_55(25)(MULT_SIZE-1) & MULT_55(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(25)(MULT_SIZE-1) & MULT_56(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(26)<=signed(MULT_55(26)(MULT_SIZE-1) & MULT_55(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(26)(MULT_SIZE-1) & MULT_56(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(27)<=signed(MULT_55(27)(MULT_SIZE-1) & MULT_55(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(27)(MULT_SIZE-1) & MULT_56(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(28)<=signed(MULT_55(28)(MULT_SIZE-1) & MULT_55(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(28)(MULT_SIZE-1) & MULT_56(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(29)<=signed(MULT_55(29)(MULT_SIZE-1) & MULT_55(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(29)(MULT_SIZE-1) & MULT_56(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(30)<=signed(MULT_55(30)(MULT_SIZE-1) & MULT_55(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(30)(MULT_SIZE-1) & MULT_56(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(31)<=signed(MULT_55(31)(MULT_SIZE-1) & MULT_55(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(31)(MULT_SIZE-1) & MULT_56(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(32)<=signed(MULT_55(32)(MULT_SIZE-1) & MULT_55(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(32)(MULT_SIZE-1) & MULT_56(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(33)<=signed(MULT_55(33)(MULT_SIZE-1) & MULT_55(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(33)(MULT_SIZE-1) & MULT_56(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(34)<=signed(MULT_55(34)(MULT_SIZE-1) & MULT_55(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(34)(MULT_SIZE-1) & MULT_56(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(35)<=signed(MULT_55(35)(MULT_SIZE-1) & MULT_55(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(35)(MULT_SIZE-1) & MULT_56(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(36)<=signed(MULT_55(36)(MULT_SIZE-1) & MULT_55(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(36)(MULT_SIZE-1) & MULT_56(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(37)<=signed(MULT_55(37)(MULT_SIZE-1) & MULT_55(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(37)(MULT_SIZE-1) & MULT_56(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(38)<=signed(MULT_55(38)(MULT_SIZE-1) & MULT_55(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(38)(MULT_SIZE-1) & MULT_56(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(39)<=signed(MULT_55(39)(MULT_SIZE-1) & MULT_55(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(39)(MULT_SIZE-1) & MULT_56(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(40)<=signed(MULT_55(40)(MULT_SIZE-1) & MULT_55(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(40)(MULT_SIZE-1) & MULT_56(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(41)<=signed(MULT_55(41)(MULT_SIZE-1) & MULT_55(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(41)(MULT_SIZE-1) & MULT_56(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(42)<=signed(MULT_55(42)(MULT_SIZE-1) & MULT_55(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(42)(MULT_SIZE-1) & MULT_56(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(43)<=signed(MULT_55(43)(MULT_SIZE-1) & MULT_55(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(43)(MULT_SIZE-1) & MULT_56(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(44)<=signed(MULT_55(44)(MULT_SIZE-1) & MULT_55(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(44)(MULT_SIZE-1) & MULT_56(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(45)<=signed(MULT_55(45)(MULT_SIZE-1) & MULT_55(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(45)(MULT_SIZE-1) & MULT_56(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(46)<=signed(MULT_55(46)(MULT_SIZE-1) & MULT_55(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(46)(MULT_SIZE-1) & MULT_56(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(47)<=signed(MULT_55(47)(MULT_SIZE-1) & MULT_55(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(47)(MULT_SIZE-1) & MULT_56(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(48)<=signed(MULT_55(48)(MULT_SIZE-1) & MULT_55(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(48)(MULT_SIZE-1) & MULT_56(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(49)<=signed(MULT_55(49)(MULT_SIZE-1) & MULT_55(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(49)(MULT_SIZE-1) & MULT_56(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(50)<=signed(MULT_55(50)(MULT_SIZE-1) & MULT_55(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(50)(MULT_SIZE-1) & MULT_56(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(51)<=signed(MULT_55(51)(MULT_SIZE-1) & MULT_55(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(51)(MULT_SIZE-1) & MULT_56(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(52)<=signed(MULT_55(52)(MULT_SIZE-1) & MULT_55(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(52)(MULT_SIZE-1) & MULT_56(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(53)<=signed(MULT_55(53)(MULT_SIZE-1) & MULT_55(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(53)(MULT_SIZE-1) & MULT_56(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(54)<=signed(MULT_55(54)(MULT_SIZE-1) & MULT_55(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(54)(MULT_SIZE-1) & MULT_56(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(55)<=signed(MULT_55(55)(MULT_SIZE-1) & MULT_55(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(55)(MULT_SIZE-1) & MULT_56(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(56)<=signed(MULT_55(56)(MULT_SIZE-1) & MULT_55(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(56)(MULT_SIZE-1) & MULT_56(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(57)<=signed(MULT_55(57)(MULT_SIZE-1) & MULT_55(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(57)(MULT_SIZE-1) & MULT_56(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(58)<=signed(MULT_55(58)(MULT_SIZE-1) & MULT_55(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(58)(MULT_SIZE-1) & MULT_56(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(59)<=signed(MULT_55(59)(MULT_SIZE-1) & MULT_55(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(59)(MULT_SIZE-1) & MULT_56(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(60)<=signed(MULT_55(60)(MULT_SIZE-1) & MULT_55(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(60)(MULT_SIZE-1) & MULT_56(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(61)<=signed(MULT_55(61)(MULT_SIZE-1) & MULT_55(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(61)(MULT_SIZE-1) & MULT_56(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(62)<=signed(MULT_55(62)(MULT_SIZE-1) & MULT_55(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(62)(MULT_SIZE-1) & MULT_56(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(63)<=signed(MULT_55(63)(MULT_SIZE-1) & MULT_55(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(63)(MULT_SIZE-1) & MULT_56(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(64)<=signed(MULT_55(64)(MULT_SIZE-1) & MULT_55(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(64)(MULT_SIZE-1) & MULT_56(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(65)<=signed(MULT_55(65)(MULT_SIZE-1) & MULT_55(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(65)(MULT_SIZE-1) & MULT_56(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(66)<=signed(MULT_55(66)(MULT_SIZE-1) & MULT_55(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(66)(MULT_SIZE-1) & MULT_56(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(67)<=signed(MULT_55(67)(MULT_SIZE-1) & MULT_55(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(67)(MULT_SIZE-1) & MULT_56(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(68)<=signed(MULT_55(68)(MULT_SIZE-1) & MULT_55(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(68)(MULT_SIZE-1) & MULT_56(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(69)<=signed(MULT_55(69)(MULT_SIZE-1) & MULT_55(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(69)(MULT_SIZE-1) & MULT_56(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(70)<=signed(MULT_55(70)(MULT_SIZE-1) & MULT_55(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(70)(MULT_SIZE-1) & MULT_56(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(71)<=signed(MULT_55(71)(MULT_SIZE-1) & MULT_55(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(71)(MULT_SIZE-1) & MULT_56(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(72)<=signed(MULT_55(72)(MULT_SIZE-1) & MULT_55(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(72)(MULT_SIZE-1) & MULT_56(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(73)<=signed(MULT_55(73)(MULT_SIZE-1) & MULT_55(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(73)(MULT_SIZE-1) & MULT_56(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(74)<=signed(MULT_55(74)(MULT_SIZE-1) & MULT_55(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(74)(MULT_SIZE-1) & MULT_56(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(75)<=signed(MULT_55(75)(MULT_SIZE-1) & MULT_55(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(75)(MULT_SIZE-1) & MULT_56(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(76)<=signed(MULT_55(76)(MULT_SIZE-1) & MULT_55(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(76)(MULT_SIZE-1) & MULT_56(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(77)<=signed(MULT_55(77)(MULT_SIZE-1) & MULT_55(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(77)(MULT_SIZE-1) & MULT_56(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(78)<=signed(MULT_55(78)(MULT_SIZE-1) & MULT_55(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(78)(MULT_SIZE-1) & MULT_56(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(79)<=signed(MULT_55(79)(MULT_SIZE-1) & MULT_55(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(79)(MULT_SIZE-1) & MULT_56(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(80)<=signed(MULT_55(80)(MULT_SIZE-1) & MULT_55(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(80)(MULT_SIZE-1) & MULT_56(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(81)<=signed(MULT_55(81)(MULT_SIZE-1) & MULT_55(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(81)(MULT_SIZE-1) & MULT_56(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(82)<=signed(MULT_55(82)(MULT_SIZE-1) & MULT_55(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(82)(MULT_SIZE-1) & MULT_56(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_28(83)<=signed(MULT_55(83)(MULT_SIZE-1) & MULT_55(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_56(83)(MULT_SIZE-1) & MULT_56(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_29(0)<=signed(MULT_57(0)(MULT_SIZE-1) & MULT_57(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(0)(MULT_SIZE-1) & MULT_58(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(1)<=signed(MULT_57(1)(MULT_SIZE-1) & MULT_57(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(1)(MULT_SIZE-1) & MULT_58(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(2)<=signed(MULT_57(2)(MULT_SIZE-1) & MULT_57(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(2)(MULT_SIZE-1) & MULT_58(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(3)<=signed(MULT_57(3)(MULT_SIZE-1) & MULT_57(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(3)(MULT_SIZE-1) & MULT_58(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(4)<=signed(MULT_57(4)(MULT_SIZE-1) & MULT_57(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(4)(MULT_SIZE-1) & MULT_58(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(5)<=signed(MULT_57(5)(MULT_SIZE-1) & MULT_57(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(5)(MULT_SIZE-1) & MULT_58(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(6)<=signed(MULT_57(6)(MULT_SIZE-1) & MULT_57(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(6)(MULT_SIZE-1) & MULT_58(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(7)<=signed(MULT_57(7)(MULT_SIZE-1) & MULT_57(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(7)(MULT_SIZE-1) & MULT_58(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(8)<=signed(MULT_57(8)(MULT_SIZE-1) & MULT_57(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(8)(MULT_SIZE-1) & MULT_58(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(9)<=signed(MULT_57(9)(MULT_SIZE-1) & MULT_57(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(9)(MULT_SIZE-1) & MULT_58(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(10)<=signed(MULT_57(10)(MULT_SIZE-1) & MULT_57(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(10)(MULT_SIZE-1) & MULT_58(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(11)<=signed(MULT_57(11)(MULT_SIZE-1) & MULT_57(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(11)(MULT_SIZE-1) & MULT_58(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(12)<=signed(MULT_57(12)(MULT_SIZE-1) & MULT_57(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(12)(MULT_SIZE-1) & MULT_58(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(13)<=signed(MULT_57(13)(MULT_SIZE-1) & MULT_57(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(13)(MULT_SIZE-1) & MULT_58(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(14)<=signed(MULT_57(14)(MULT_SIZE-1) & MULT_57(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(14)(MULT_SIZE-1) & MULT_58(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(15)<=signed(MULT_57(15)(MULT_SIZE-1) & MULT_57(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(15)(MULT_SIZE-1) & MULT_58(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(16)<=signed(MULT_57(16)(MULT_SIZE-1) & MULT_57(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(16)(MULT_SIZE-1) & MULT_58(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(17)<=signed(MULT_57(17)(MULT_SIZE-1) & MULT_57(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(17)(MULT_SIZE-1) & MULT_58(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(18)<=signed(MULT_57(18)(MULT_SIZE-1) & MULT_57(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(18)(MULT_SIZE-1) & MULT_58(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(19)<=signed(MULT_57(19)(MULT_SIZE-1) & MULT_57(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(19)(MULT_SIZE-1) & MULT_58(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(20)<=signed(MULT_57(20)(MULT_SIZE-1) & MULT_57(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(20)(MULT_SIZE-1) & MULT_58(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(21)<=signed(MULT_57(21)(MULT_SIZE-1) & MULT_57(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(21)(MULT_SIZE-1) & MULT_58(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(22)<=signed(MULT_57(22)(MULT_SIZE-1) & MULT_57(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(22)(MULT_SIZE-1) & MULT_58(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(23)<=signed(MULT_57(23)(MULT_SIZE-1) & MULT_57(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(23)(MULT_SIZE-1) & MULT_58(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(24)<=signed(MULT_57(24)(MULT_SIZE-1) & MULT_57(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(24)(MULT_SIZE-1) & MULT_58(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(25)<=signed(MULT_57(25)(MULT_SIZE-1) & MULT_57(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(25)(MULT_SIZE-1) & MULT_58(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(26)<=signed(MULT_57(26)(MULT_SIZE-1) & MULT_57(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(26)(MULT_SIZE-1) & MULT_58(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(27)<=signed(MULT_57(27)(MULT_SIZE-1) & MULT_57(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(27)(MULT_SIZE-1) & MULT_58(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(28)<=signed(MULT_57(28)(MULT_SIZE-1) & MULT_57(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(28)(MULT_SIZE-1) & MULT_58(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(29)<=signed(MULT_57(29)(MULT_SIZE-1) & MULT_57(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(29)(MULT_SIZE-1) & MULT_58(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(30)<=signed(MULT_57(30)(MULT_SIZE-1) & MULT_57(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(30)(MULT_SIZE-1) & MULT_58(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(31)<=signed(MULT_57(31)(MULT_SIZE-1) & MULT_57(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(31)(MULT_SIZE-1) & MULT_58(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(32)<=signed(MULT_57(32)(MULT_SIZE-1) & MULT_57(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(32)(MULT_SIZE-1) & MULT_58(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(33)<=signed(MULT_57(33)(MULT_SIZE-1) & MULT_57(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(33)(MULT_SIZE-1) & MULT_58(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(34)<=signed(MULT_57(34)(MULT_SIZE-1) & MULT_57(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(34)(MULT_SIZE-1) & MULT_58(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(35)<=signed(MULT_57(35)(MULT_SIZE-1) & MULT_57(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(35)(MULT_SIZE-1) & MULT_58(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(36)<=signed(MULT_57(36)(MULT_SIZE-1) & MULT_57(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(36)(MULT_SIZE-1) & MULT_58(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(37)<=signed(MULT_57(37)(MULT_SIZE-1) & MULT_57(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(37)(MULT_SIZE-1) & MULT_58(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(38)<=signed(MULT_57(38)(MULT_SIZE-1) & MULT_57(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(38)(MULT_SIZE-1) & MULT_58(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(39)<=signed(MULT_57(39)(MULT_SIZE-1) & MULT_57(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(39)(MULT_SIZE-1) & MULT_58(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(40)<=signed(MULT_57(40)(MULT_SIZE-1) & MULT_57(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(40)(MULT_SIZE-1) & MULT_58(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(41)<=signed(MULT_57(41)(MULT_SIZE-1) & MULT_57(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(41)(MULT_SIZE-1) & MULT_58(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(42)<=signed(MULT_57(42)(MULT_SIZE-1) & MULT_57(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(42)(MULT_SIZE-1) & MULT_58(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(43)<=signed(MULT_57(43)(MULT_SIZE-1) & MULT_57(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(43)(MULT_SIZE-1) & MULT_58(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(44)<=signed(MULT_57(44)(MULT_SIZE-1) & MULT_57(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(44)(MULT_SIZE-1) & MULT_58(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(45)<=signed(MULT_57(45)(MULT_SIZE-1) & MULT_57(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(45)(MULT_SIZE-1) & MULT_58(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(46)<=signed(MULT_57(46)(MULT_SIZE-1) & MULT_57(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(46)(MULT_SIZE-1) & MULT_58(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(47)<=signed(MULT_57(47)(MULT_SIZE-1) & MULT_57(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(47)(MULT_SIZE-1) & MULT_58(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(48)<=signed(MULT_57(48)(MULT_SIZE-1) & MULT_57(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(48)(MULT_SIZE-1) & MULT_58(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(49)<=signed(MULT_57(49)(MULT_SIZE-1) & MULT_57(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(49)(MULT_SIZE-1) & MULT_58(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(50)<=signed(MULT_57(50)(MULT_SIZE-1) & MULT_57(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(50)(MULT_SIZE-1) & MULT_58(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(51)<=signed(MULT_57(51)(MULT_SIZE-1) & MULT_57(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(51)(MULT_SIZE-1) & MULT_58(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(52)<=signed(MULT_57(52)(MULT_SIZE-1) & MULT_57(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(52)(MULT_SIZE-1) & MULT_58(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(53)<=signed(MULT_57(53)(MULT_SIZE-1) & MULT_57(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(53)(MULT_SIZE-1) & MULT_58(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(54)<=signed(MULT_57(54)(MULT_SIZE-1) & MULT_57(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(54)(MULT_SIZE-1) & MULT_58(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(55)<=signed(MULT_57(55)(MULT_SIZE-1) & MULT_57(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(55)(MULT_SIZE-1) & MULT_58(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(56)<=signed(MULT_57(56)(MULT_SIZE-1) & MULT_57(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(56)(MULT_SIZE-1) & MULT_58(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(57)<=signed(MULT_57(57)(MULT_SIZE-1) & MULT_57(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(57)(MULT_SIZE-1) & MULT_58(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(58)<=signed(MULT_57(58)(MULT_SIZE-1) & MULT_57(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(58)(MULT_SIZE-1) & MULT_58(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(59)<=signed(MULT_57(59)(MULT_SIZE-1) & MULT_57(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(59)(MULT_SIZE-1) & MULT_58(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(60)<=signed(MULT_57(60)(MULT_SIZE-1) & MULT_57(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(60)(MULT_SIZE-1) & MULT_58(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(61)<=signed(MULT_57(61)(MULT_SIZE-1) & MULT_57(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(61)(MULT_SIZE-1) & MULT_58(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(62)<=signed(MULT_57(62)(MULT_SIZE-1) & MULT_57(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(62)(MULT_SIZE-1) & MULT_58(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(63)<=signed(MULT_57(63)(MULT_SIZE-1) & MULT_57(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(63)(MULT_SIZE-1) & MULT_58(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(64)<=signed(MULT_57(64)(MULT_SIZE-1) & MULT_57(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(64)(MULT_SIZE-1) & MULT_58(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(65)<=signed(MULT_57(65)(MULT_SIZE-1) & MULT_57(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(65)(MULT_SIZE-1) & MULT_58(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(66)<=signed(MULT_57(66)(MULT_SIZE-1) & MULT_57(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(66)(MULT_SIZE-1) & MULT_58(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(67)<=signed(MULT_57(67)(MULT_SIZE-1) & MULT_57(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(67)(MULT_SIZE-1) & MULT_58(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(68)<=signed(MULT_57(68)(MULT_SIZE-1) & MULT_57(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(68)(MULT_SIZE-1) & MULT_58(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(69)<=signed(MULT_57(69)(MULT_SIZE-1) & MULT_57(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(69)(MULT_SIZE-1) & MULT_58(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(70)<=signed(MULT_57(70)(MULT_SIZE-1) & MULT_57(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(70)(MULT_SIZE-1) & MULT_58(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(71)<=signed(MULT_57(71)(MULT_SIZE-1) & MULT_57(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(71)(MULT_SIZE-1) & MULT_58(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(72)<=signed(MULT_57(72)(MULT_SIZE-1) & MULT_57(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(72)(MULT_SIZE-1) & MULT_58(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(73)<=signed(MULT_57(73)(MULT_SIZE-1) & MULT_57(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(73)(MULT_SIZE-1) & MULT_58(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(74)<=signed(MULT_57(74)(MULT_SIZE-1) & MULT_57(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(74)(MULT_SIZE-1) & MULT_58(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(75)<=signed(MULT_57(75)(MULT_SIZE-1) & MULT_57(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(75)(MULT_SIZE-1) & MULT_58(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(76)<=signed(MULT_57(76)(MULT_SIZE-1) & MULT_57(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(76)(MULT_SIZE-1) & MULT_58(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(77)<=signed(MULT_57(77)(MULT_SIZE-1) & MULT_57(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(77)(MULT_SIZE-1) & MULT_58(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(78)<=signed(MULT_57(78)(MULT_SIZE-1) & MULT_57(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(78)(MULT_SIZE-1) & MULT_58(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(79)<=signed(MULT_57(79)(MULT_SIZE-1) & MULT_57(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(79)(MULT_SIZE-1) & MULT_58(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(80)<=signed(MULT_57(80)(MULT_SIZE-1) & MULT_57(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(80)(MULT_SIZE-1) & MULT_58(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(81)<=signed(MULT_57(81)(MULT_SIZE-1) & MULT_57(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(81)(MULT_SIZE-1) & MULT_58(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(82)<=signed(MULT_57(82)(MULT_SIZE-1) & MULT_57(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(82)(MULT_SIZE-1) & MULT_58(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_29(83)<=signed(MULT_57(83)(MULT_SIZE-1) & MULT_57(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_58(83)(MULT_SIZE-1) & MULT_58(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_30(0)<=signed(MULT_59(0)(MULT_SIZE-1) & MULT_59(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(0)(MULT_SIZE-1) & MULT_60(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(1)<=signed(MULT_59(1)(MULT_SIZE-1) & MULT_59(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(1)(MULT_SIZE-1) & MULT_60(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(2)<=signed(MULT_59(2)(MULT_SIZE-1) & MULT_59(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(2)(MULT_SIZE-1) & MULT_60(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(3)<=signed(MULT_59(3)(MULT_SIZE-1) & MULT_59(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(3)(MULT_SIZE-1) & MULT_60(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(4)<=signed(MULT_59(4)(MULT_SIZE-1) & MULT_59(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(4)(MULT_SIZE-1) & MULT_60(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(5)<=signed(MULT_59(5)(MULT_SIZE-1) & MULT_59(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(5)(MULT_SIZE-1) & MULT_60(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(6)<=signed(MULT_59(6)(MULT_SIZE-1) & MULT_59(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(6)(MULT_SIZE-1) & MULT_60(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(7)<=signed(MULT_59(7)(MULT_SIZE-1) & MULT_59(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(7)(MULT_SIZE-1) & MULT_60(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(8)<=signed(MULT_59(8)(MULT_SIZE-1) & MULT_59(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(8)(MULT_SIZE-1) & MULT_60(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(9)<=signed(MULT_59(9)(MULT_SIZE-1) & MULT_59(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(9)(MULT_SIZE-1) & MULT_60(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(10)<=signed(MULT_59(10)(MULT_SIZE-1) & MULT_59(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(10)(MULT_SIZE-1) & MULT_60(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(11)<=signed(MULT_59(11)(MULT_SIZE-1) & MULT_59(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(11)(MULT_SIZE-1) & MULT_60(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(12)<=signed(MULT_59(12)(MULT_SIZE-1) & MULT_59(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(12)(MULT_SIZE-1) & MULT_60(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(13)<=signed(MULT_59(13)(MULT_SIZE-1) & MULT_59(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(13)(MULT_SIZE-1) & MULT_60(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(14)<=signed(MULT_59(14)(MULT_SIZE-1) & MULT_59(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(14)(MULT_SIZE-1) & MULT_60(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(15)<=signed(MULT_59(15)(MULT_SIZE-1) & MULT_59(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(15)(MULT_SIZE-1) & MULT_60(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(16)<=signed(MULT_59(16)(MULT_SIZE-1) & MULT_59(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(16)(MULT_SIZE-1) & MULT_60(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(17)<=signed(MULT_59(17)(MULT_SIZE-1) & MULT_59(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(17)(MULT_SIZE-1) & MULT_60(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(18)<=signed(MULT_59(18)(MULT_SIZE-1) & MULT_59(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(18)(MULT_SIZE-1) & MULT_60(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(19)<=signed(MULT_59(19)(MULT_SIZE-1) & MULT_59(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(19)(MULT_SIZE-1) & MULT_60(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(20)<=signed(MULT_59(20)(MULT_SIZE-1) & MULT_59(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(20)(MULT_SIZE-1) & MULT_60(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(21)<=signed(MULT_59(21)(MULT_SIZE-1) & MULT_59(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(21)(MULT_SIZE-1) & MULT_60(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(22)<=signed(MULT_59(22)(MULT_SIZE-1) & MULT_59(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(22)(MULT_SIZE-1) & MULT_60(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(23)<=signed(MULT_59(23)(MULT_SIZE-1) & MULT_59(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(23)(MULT_SIZE-1) & MULT_60(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(24)<=signed(MULT_59(24)(MULT_SIZE-1) & MULT_59(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(24)(MULT_SIZE-1) & MULT_60(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(25)<=signed(MULT_59(25)(MULT_SIZE-1) & MULT_59(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(25)(MULT_SIZE-1) & MULT_60(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(26)<=signed(MULT_59(26)(MULT_SIZE-1) & MULT_59(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(26)(MULT_SIZE-1) & MULT_60(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(27)<=signed(MULT_59(27)(MULT_SIZE-1) & MULT_59(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(27)(MULT_SIZE-1) & MULT_60(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(28)<=signed(MULT_59(28)(MULT_SIZE-1) & MULT_59(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(28)(MULT_SIZE-1) & MULT_60(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(29)<=signed(MULT_59(29)(MULT_SIZE-1) & MULT_59(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(29)(MULT_SIZE-1) & MULT_60(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(30)<=signed(MULT_59(30)(MULT_SIZE-1) & MULT_59(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(30)(MULT_SIZE-1) & MULT_60(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(31)<=signed(MULT_59(31)(MULT_SIZE-1) & MULT_59(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(31)(MULT_SIZE-1) & MULT_60(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(32)<=signed(MULT_59(32)(MULT_SIZE-1) & MULT_59(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(32)(MULT_SIZE-1) & MULT_60(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(33)<=signed(MULT_59(33)(MULT_SIZE-1) & MULT_59(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(33)(MULT_SIZE-1) & MULT_60(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(34)<=signed(MULT_59(34)(MULT_SIZE-1) & MULT_59(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(34)(MULT_SIZE-1) & MULT_60(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(35)<=signed(MULT_59(35)(MULT_SIZE-1) & MULT_59(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(35)(MULT_SIZE-1) & MULT_60(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(36)<=signed(MULT_59(36)(MULT_SIZE-1) & MULT_59(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(36)(MULT_SIZE-1) & MULT_60(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(37)<=signed(MULT_59(37)(MULT_SIZE-1) & MULT_59(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(37)(MULT_SIZE-1) & MULT_60(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(38)<=signed(MULT_59(38)(MULT_SIZE-1) & MULT_59(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(38)(MULT_SIZE-1) & MULT_60(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(39)<=signed(MULT_59(39)(MULT_SIZE-1) & MULT_59(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(39)(MULT_SIZE-1) & MULT_60(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(40)<=signed(MULT_59(40)(MULT_SIZE-1) & MULT_59(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(40)(MULT_SIZE-1) & MULT_60(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(41)<=signed(MULT_59(41)(MULT_SIZE-1) & MULT_59(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(41)(MULT_SIZE-1) & MULT_60(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(42)<=signed(MULT_59(42)(MULT_SIZE-1) & MULT_59(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(42)(MULT_SIZE-1) & MULT_60(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(43)<=signed(MULT_59(43)(MULT_SIZE-1) & MULT_59(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(43)(MULT_SIZE-1) & MULT_60(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(44)<=signed(MULT_59(44)(MULT_SIZE-1) & MULT_59(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(44)(MULT_SIZE-1) & MULT_60(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(45)<=signed(MULT_59(45)(MULT_SIZE-1) & MULT_59(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(45)(MULT_SIZE-1) & MULT_60(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(46)<=signed(MULT_59(46)(MULT_SIZE-1) & MULT_59(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(46)(MULT_SIZE-1) & MULT_60(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(47)<=signed(MULT_59(47)(MULT_SIZE-1) & MULT_59(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(47)(MULT_SIZE-1) & MULT_60(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(48)<=signed(MULT_59(48)(MULT_SIZE-1) & MULT_59(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(48)(MULT_SIZE-1) & MULT_60(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(49)<=signed(MULT_59(49)(MULT_SIZE-1) & MULT_59(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(49)(MULT_SIZE-1) & MULT_60(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(50)<=signed(MULT_59(50)(MULT_SIZE-1) & MULT_59(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(50)(MULT_SIZE-1) & MULT_60(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(51)<=signed(MULT_59(51)(MULT_SIZE-1) & MULT_59(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(51)(MULT_SIZE-1) & MULT_60(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(52)<=signed(MULT_59(52)(MULT_SIZE-1) & MULT_59(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(52)(MULT_SIZE-1) & MULT_60(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(53)<=signed(MULT_59(53)(MULT_SIZE-1) & MULT_59(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(53)(MULT_SIZE-1) & MULT_60(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(54)<=signed(MULT_59(54)(MULT_SIZE-1) & MULT_59(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(54)(MULT_SIZE-1) & MULT_60(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(55)<=signed(MULT_59(55)(MULT_SIZE-1) & MULT_59(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(55)(MULT_SIZE-1) & MULT_60(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(56)<=signed(MULT_59(56)(MULT_SIZE-1) & MULT_59(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(56)(MULT_SIZE-1) & MULT_60(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(57)<=signed(MULT_59(57)(MULT_SIZE-1) & MULT_59(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(57)(MULT_SIZE-1) & MULT_60(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(58)<=signed(MULT_59(58)(MULT_SIZE-1) & MULT_59(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(58)(MULT_SIZE-1) & MULT_60(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(59)<=signed(MULT_59(59)(MULT_SIZE-1) & MULT_59(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(59)(MULT_SIZE-1) & MULT_60(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(60)<=signed(MULT_59(60)(MULT_SIZE-1) & MULT_59(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(60)(MULT_SIZE-1) & MULT_60(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(61)<=signed(MULT_59(61)(MULT_SIZE-1) & MULT_59(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(61)(MULT_SIZE-1) & MULT_60(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(62)<=signed(MULT_59(62)(MULT_SIZE-1) & MULT_59(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(62)(MULT_SIZE-1) & MULT_60(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(63)<=signed(MULT_59(63)(MULT_SIZE-1) & MULT_59(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(63)(MULT_SIZE-1) & MULT_60(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(64)<=signed(MULT_59(64)(MULT_SIZE-1) & MULT_59(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(64)(MULT_SIZE-1) & MULT_60(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(65)<=signed(MULT_59(65)(MULT_SIZE-1) & MULT_59(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(65)(MULT_SIZE-1) & MULT_60(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(66)<=signed(MULT_59(66)(MULT_SIZE-1) & MULT_59(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(66)(MULT_SIZE-1) & MULT_60(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(67)<=signed(MULT_59(67)(MULT_SIZE-1) & MULT_59(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(67)(MULT_SIZE-1) & MULT_60(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(68)<=signed(MULT_59(68)(MULT_SIZE-1) & MULT_59(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(68)(MULT_SIZE-1) & MULT_60(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(69)<=signed(MULT_59(69)(MULT_SIZE-1) & MULT_59(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(69)(MULT_SIZE-1) & MULT_60(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(70)<=signed(MULT_59(70)(MULT_SIZE-1) & MULT_59(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(70)(MULT_SIZE-1) & MULT_60(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(71)<=signed(MULT_59(71)(MULT_SIZE-1) & MULT_59(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(71)(MULT_SIZE-1) & MULT_60(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(72)<=signed(MULT_59(72)(MULT_SIZE-1) & MULT_59(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(72)(MULT_SIZE-1) & MULT_60(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(73)<=signed(MULT_59(73)(MULT_SIZE-1) & MULT_59(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(73)(MULT_SIZE-1) & MULT_60(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(74)<=signed(MULT_59(74)(MULT_SIZE-1) & MULT_59(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(74)(MULT_SIZE-1) & MULT_60(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(75)<=signed(MULT_59(75)(MULT_SIZE-1) & MULT_59(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(75)(MULT_SIZE-1) & MULT_60(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(76)<=signed(MULT_59(76)(MULT_SIZE-1) & MULT_59(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(76)(MULT_SIZE-1) & MULT_60(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(77)<=signed(MULT_59(77)(MULT_SIZE-1) & MULT_59(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(77)(MULT_SIZE-1) & MULT_60(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(78)<=signed(MULT_59(78)(MULT_SIZE-1) & MULT_59(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(78)(MULT_SIZE-1) & MULT_60(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(79)<=signed(MULT_59(79)(MULT_SIZE-1) & MULT_59(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(79)(MULT_SIZE-1) & MULT_60(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(80)<=signed(MULT_59(80)(MULT_SIZE-1) & MULT_59(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(80)(MULT_SIZE-1) & MULT_60(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(81)<=signed(MULT_59(81)(MULT_SIZE-1) & MULT_59(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(81)(MULT_SIZE-1) & MULT_60(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(82)<=signed(MULT_59(82)(MULT_SIZE-1) & MULT_59(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(82)(MULT_SIZE-1) & MULT_60(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_30(83)<=signed(MULT_59(83)(MULT_SIZE-1) & MULT_59(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_60(83)(MULT_SIZE-1) & MULT_60(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_31(0)<=signed(MULT_61(0)(MULT_SIZE-1) & MULT_61(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(0)(MULT_SIZE-1) & MULT_62(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(1)<=signed(MULT_61(1)(MULT_SIZE-1) & MULT_61(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(1)(MULT_SIZE-1) & MULT_62(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(2)<=signed(MULT_61(2)(MULT_SIZE-1) & MULT_61(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(2)(MULT_SIZE-1) & MULT_62(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(3)<=signed(MULT_61(3)(MULT_SIZE-1) & MULT_61(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(3)(MULT_SIZE-1) & MULT_62(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(4)<=signed(MULT_61(4)(MULT_SIZE-1) & MULT_61(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(4)(MULT_SIZE-1) & MULT_62(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(5)<=signed(MULT_61(5)(MULT_SIZE-1) & MULT_61(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(5)(MULT_SIZE-1) & MULT_62(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(6)<=signed(MULT_61(6)(MULT_SIZE-1) & MULT_61(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(6)(MULT_SIZE-1) & MULT_62(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(7)<=signed(MULT_61(7)(MULT_SIZE-1) & MULT_61(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(7)(MULT_SIZE-1) & MULT_62(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(8)<=signed(MULT_61(8)(MULT_SIZE-1) & MULT_61(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(8)(MULT_SIZE-1) & MULT_62(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(9)<=signed(MULT_61(9)(MULT_SIZE-1) & MULT_61(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(9)(MULT_SIZE-1) & MULT_62(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(10)<=signed(MULT_61(10)(MULT_SIZE-1) & MULT_61(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(10)(MULT_SIZE-1) & MULT_62(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(11)<=signed(MULT_61(11)(MULT_SIZE-1) & MULT_61(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(11)(MULT_SIZE-1) & MULT_62(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(12)<=signed(MULT_61(12)(MULT_SIZE-1) & MULT_61(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(12)(MULT_SIZE-1) & MULT_62(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(13)<=signed(MULT_61(13)(MULT_SIZE-1) & MULT_61(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(13)(MULT_SIZE-1) & MULT_62(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(14)<=signed(MULT_61(14)(MULT_SIZE-1) & MULT_61(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(14)(MULT_SIZE-1) & MULT_62(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(15)<=signed(MULT_61(15)(MULT_SIZE-1) & MULT_61(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(15)(MULT_SIZE-1) & MULT_62(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(16)<=signed(MULT_61(16)(MULT_SIZE-1) & MULT_61(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(16)(MULT_SIZE-1) & MULT_62(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(17)<=signed(MULT_61(17)(MULT_SIZE-1) & MULT_61(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(17)(MULT_SIZE-1) & MULT_62(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(18)<=signed(MULT_61(18)(MULT_SIZE-1) & MULT_61(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(18)(MULT_SIZE-1) & MULT_62(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(19)<=signed(MULT_61(19)(MULT_SIZE-1) & MULT_61(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(19)(MULT_SIZE-1) & MULT_62(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(20)<=signed(MULT_61(20)(MULT_SIZE-1) & MULT_61(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(20)(MULT_SIZE-1) & MULT_62(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(21)<=signed(MULT_61(21)(MULT_SIZE-1) & MULT_61(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(21)(MULT_SIZE-1) & MULT_62(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(22)<=signed(MULT_61(22)(MULT_SIZE-1) & MULT_61(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(22)(MULT_SIZE-1) & MULT_62(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(23)<=signed(MULT_61(23)(MULT_SIZE-1) & MULT_61(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(23)(MULT_SIZE-1) & MULT_62(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(24)<=signed(MULT_61(24)(MULT_SIZE-1) & MULT_61(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(24)(MULT_SIZE-1) & MULT_62(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(25)<=signed(MULT_61(25)(MULT_SIZE-1) & MULT_61(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(25)(MULT_SIZE-1) & MULT_62(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(26)<=signed(MULT_61(26)(MULT_SIZE-1) & MULT_61(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(26)(MULT_SIZE-1) & MULT_62(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(27)<=signed(MULT_61(27)(MULT_SIZE-1) & MULT_61(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(27)(MULT_SIZE-1) & MULT_62(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(28)<=signed(MULT_61(28)(MULT_SIZE-1) & MULT_61(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(28)(MULT_SIZE-1) & MULT_62(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(29)<=signed(MULT_61(29)(MULT_SIZE-1) & MULT_61(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(29)(MULT_SIZE-1) & MULT_62(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(30)<=signed(MULT_61(30)(MULT_SIZE-1) & MULT_61(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(30)(MULT_SIZE-1) & MULT_62(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(31)<=signed(MULT_61(31)(MULT_SIZE-1) & MULT_61(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(31)(MULT_SIZE-1) & MULT_62(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(32)<=signed(MULT_61(32)(MULT_SIZE-1) & MULT_61(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(32)(MULT_SIZE-1) & MULT_62(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(33)<=signed(MULT_61(33)(MULT_SIZE-1) & MULT_61(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(33)(MULT_SIZE-1) & MULT_62(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(34)<=signed(MULT_61(34)(MULT_SIZE-1) & MULT_61(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(34)(MULT_SIZE-1) & MULT_62(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(35)<=signed(MULT_61(35)(MULT_SIZE-1) & MULT_61(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(35)(MULT_SIZE-1) & MULT_62(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(36)<=signed(MULT_61(36)(MULT_SIZE-1) & MULT_61(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(36)(MULT_SIZE-1) & MULT_62(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(37)<=signed(MULT_61(37)(MULT_SIZE-1) & MULT_61(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(37)(MULT_SIZE-1) & MULT_62(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(38)<=signed(MULT_61(38)(MULT_SIZE-1) & MULT_61(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(38)(MULT_SIZE-1) & MULT_62(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(39)<=signed(MULT_61(39)(MULT_SIZE-1) & MULT_61(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(39)(MULT_SIZE-1) & MULT_62(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(40)<=signed(MULT_61(40)(MULT_SIZE-1) & MULT_61(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(40)(MULT_SIZE-1) & MULT_62(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(41)<=signed(MULT_61(41)(MULT_SIZE-1) & MULT_61(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(41)(MULT_SIZE-1) & MULT_62(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(42)<=signed(MULT_61(42)(MULT_SIZE-1) & MULT_61(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(42)(MULT_SIZE-1) & MULT_62(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(43)<=signed(MULT_61(43)(MULT_SIZE-1) & MULT_61(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(43)(MULT_SIZE-1) & MULT_62(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(44)<=signed(MULT_61(44)(MULT_SIZE-1) & MULT_61(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(44)(MULT_SIZE-1) & MULT_62(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(45)<=signed(MULT_61(45)(MULT_SIZE-1) & MULT_61(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(45)(MULT_SIZE-1) & MULT_62(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(46)<=signed(MULT_61(46)(MULT_SIZE-1) & MULT_61(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(46)(MULT_SIZE-1) & MULT_62(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(47)<=signed(MULT_61(47)(MULT_SIZE-1) & MULT_61(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(47)(MULT_SIZE-1) & MULT_62(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(48)<=signed(MULT_61(48)(MULT_SIZE-1) & MULT_61(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(48)(MULT_SIZE-1) & MULT_62(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(49)<=signed(MULT_61(49)(MULT_SIZE-1) & MULT_61(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(49)(MULT_SIZE-1) & MULT_62(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(50)<=signed(MULT_61(50)(MULT_SIZE-1) & MULT_61(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(50)(MULT_SIZE-1) & MULT_62(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(51)<=signed(MULT_61(51)(MULT_SIZE-1) & MULT_61(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(51)(MULT_SIZE-1) & MULT_62(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(52)<=signed(MULT_61(52)(MULT_SIZE-1) & MULT_61(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(52)(MULT_SIZE-1) & MULT_62(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(53)<=signed(MULT_61(53)(MULT_SIZE-1) & MULT_61(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(53)(MULT_SIZE-1) & MULT_62(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(54)<=signed(MULT_61(54)(MULT_SIZE-1) & MULT_61(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(54)(MULT_SIZE-1) & MULT_62(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(55)<=signed(MULT_61(55)(MULT_SIZE-1) & MULT_61(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(55)(MULT_SIZE-1) & MULT_62(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(56)<=signed(MULT_61(56)(MULT_SIZE-1) & MULT_61(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(56)(MULT_SIZE-1) & MULT_62(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(57)<=signed(MULT_61(57)(MULT_SIZE-1) & MULT_61(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(57)(MULT_SIZE-1) & MULT_62(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(58)<=signed(MULT_61(58)(MULT_SIZE-1) & MULT_61(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(58)(MULT_SIZE-1) & MULT_62(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(59)<=signed(MULT_61(59)(MULT_SIZE-1) & MULT_61(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(59)(MULT_SIZE-1) & MULT_62(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(60)<=signed(MULT_61(60)(MULT_SIZE-1) & MULT_61(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(60)(MULT_SIZE-1) & MULT_62(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(61)<=signed(MULT_61(61)(MULT_SIZE-1) & MULT_61(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(61)(MULT_SIZE-1) & MULT_62(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(62)<=signed(MULT_61(62)(MULT_SIZE-1) & MULT_61(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(62)(MULT_SIZE-1) & MULT_62(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(63)<=signed(MULT_61(63)(MULT_SIZE-1) & MULT_61(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(63)(MULT_SIZE-1) & MULT_62(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(64)<=signed(MULT_61(64)(MULT_SIZE-1) & MULT_61(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(64)(MULT_SIZE-1) & MULT_62(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(65)<=signed(MULT_61(65)(MULT_SIZE-1) & MULT_61(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(65)(MULT_SIZE-1) & MULT_62(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(66)<=signed(MULT_61(66)(MULT_SIZE-1) & MULT_61(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(66)(MULT_SIZE-1) & MULT_62(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(67)<=signed(MULT_61(67)(MULT_SIZE-1) & MULT_61(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(67)(MULT_SIZE-1) & MULT_62(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(68)<=signed(MULT_61(68)(MULT_SIZE-1) & MULT_61(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(68)(MULT_SIZE-1) & MULT_62(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(69)<=signed(MULT_61(69)(MULT_SIZE-1) & MULT_61(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(69)(MULT_SIZE-1) & MULT_62(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(70)<=signed(MULT_61(70)(MULT_SIZE-1) & MULT_61(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(70)(MULT_SIZE-1) & MULT_62(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(71)<=signed(MULT_61(71)(MULT_SIZE-1) & MULT_61(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(71)(MULT_SIZE-1) & MULT_62(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(72)<=signed(MULT_61(72)(MULT_SIZE-1) & MULT_61(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(72)(MULT_SIZE-1) & MULT_62(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(73)<=signed(MULT_61(73)(MULT_SIZE-1) & MULT_61(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(73)(MULT_SIZE-1) & MULT_62(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(74)<=signed(MULT_61(74)(MULT_SIZE-1) & MULT_61(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(74)(MULT_SIZE-1) & MULT_62(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(75)<=signed(MULT_61(75)(MULT_SIZE-1) & MULT_61(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(75)(MULT_SIZE-1) & MULT_62(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(76)<=signed(MULT_61(76)(MULT_SIZE-1) & MULT_61(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(76)(MULT_SIZE-1) & MULT_62(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(77)<=signed(MULT_61(77)(MULT_SIZE-1) & MULT_61(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(77)(MULT_SIZE-1) & MULT_62(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(78)<=signed(MULT_61(78)(MULT_SIZE-1) & MULT_61(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(78)(MULT_SIZE-1) & MULT_62(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(79)<=signed(MULT_61(79)(MULT_SIZE-1) & MULT_61(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(79)(MULT_SIZE-1) & MULT_62(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(80)<=signed(MULT_61(80)(MULT_SIZE-1) & MULT_61(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(80)(MULT_SIZE-1) & MULT_62(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(81)<=signed(MULT_61(81)(MULT_SIZE-1) & MULT_61(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(81)(MULT_SIZE-1) & MULT_62(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(82)<=signed(MULT_61(82)(MULT_SIZE-1) & MULT_61(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(82)(MULT_SIZE-1) & MULT_62(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_31(83)<=signed(MULT_61(83)(MULT_SIZE-1) & MULT_61(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_62(83)(MULT_SIZE-1) & MULT_62(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_32(0)<=signed(MULT_63(0)(MULT_SIZE-1) & MULT_63(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(0)(MULT_SIZE-1) & MULT_64(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(1)<=signed(MULT_63(1)(MULT_SIZE-1) & MULT_63(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(1)(MULT_SIZE-1) & MULT_64(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(2)<=signed(MULT_63(2)(MULT_SIZE-1) & MULT_63(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(2)(MULT_SIZE-1) & MULT_64(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(3)<=signed(MULT_63(3)(MULT_SIZE-1) & MULT_63(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(3)(MULT_SIZE-1) & MULT_64(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(4)<=signed(MULT_63(4)(MULT_SIZE-1) & MULT_63(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(4)(MULT_SIZE-1) & MULT_64(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(5)<=signed(MULT_63(5)(MULT_SIZE-1) & MULT_63(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(5)(MULT_SIZE-1) & MULT_64(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(6)<=signed(MULT_63(6)(MULT_SIZE-1) & MULT_63(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(6)(MULT_SIZE-1) & MULT_64(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(7)<=signed(MULT_63(7)(MULT_SIZE-1) & MULT_63(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(7)(MULT_SIZE-1) & MULT_64(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(8)<=signed(MULT_63(8)(MULT_SIZE-1) & MULT_63(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(8)(MULT_SIZE-1) & MULT_64(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(9)<=signed(MULT_63(9)(MULT_SIZE-1) & MULT_63(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(9)(MULT_SIZE-1) & MULT_64(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(10)<=signed(MULT_63(10)(MULT_SIZE-1) & MULT_63(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(10)(MULT_SIZE-1) & MULT_64(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(11)<=signed(MULT_63(11)(MULT_SIZE-1) & MULT_63(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(11)(MULT_SIZE-1) & MULT_64(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(12)<=signed(MULT_63(12)(MULT_SIZE-1) & MULT_63(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(12)(MULT_SIZE-1) & MULT_64(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(13)<=signed(MULT_63(13)(MULT_SIZE-1) & MULT_63(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(13)(MULT_SIZE-1) & MULT_64(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(14)<=signed(MULT_63(14)(MULT_SIZE-1) & MULT_63(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(14)(MULT_SIZE-1) & MULT_64(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(15)<=signed(MULT_63(15)(MULT_SIZE-1) & MULT_63(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(15)(MULT_SIZE-1) & MULT_64(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(16)<=signed(MULT_63(16)(MULT_SIZE-1) & MULT_63(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(16)(MULT_SIZE-1) & MULT_64(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(17)<=signed(MULT_63(17)(MULT_SIZE-1) & MULT_63(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(17)(MULT_SIZE-1) & MULT_64(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(18)<=signed(MULT_63(18)(MULT_SIZE-1) & MULT_63(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(18)(MULT_SIZE-1) & MULT_64(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(19)<=signed(MULT_63(19)(MULT_SIZE-1) & MULT_63(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(19)(MULT_SIZE-1) & MULT_64(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(20)<=signed(MULT_63(20)(MULT_SIZE-1) & MULT_63(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(20)(MULT_SIZE-1) & MULT_64(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(21)<=signed(MULT_63(21)(MULT_SIZE-1) & MULT_63(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(21)(MULT_SIZE-1) & MULT_64(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(22)<=signed(MULT_63(22)(MULT_SIZE-1) & MULT_63(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(22)(MULT_SIZE-1) & MULT_64(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(23)<=signed(MULT_63(23)(MULT_SIZE-1) & MULT_63(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(23)(MULT_SIZE-1) & MULT_64(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(24)<=signed(MULT_63(24)(MULT_SIZE-1) & MULT_63(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(24)(MULT_SIZE-1) & MULT_64(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(25)<=signed(MULT_63(25)(MULT_SIZE-1) & MULT_63(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(25)(MULT_SIZE-1) & MULT_64(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(26)<=signed(MULT_63(26)(MULT_SIZE-1) & MULT_63(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(26)(MULT_SIZE-1) & MULT_64(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(27)<=signed(MULT_63(27)(MULT_SIZE-1) & MULT_63(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(27)(MULT_SIZE-1) & MULT_64(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(28)<=signed(MULT_63(28)(MULT_SIZE-1) & MULT_63(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(28)(MULT_SIZE-1) & MULT_64(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(29)<=signed(MULT_63(29)(MULT_SIZE-1) & MULT_63(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(29)(MULT_SIZE-1) & MULT_64(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(30)<=signed(MULT_63(30)(MULT_SIZE-1) & MULT_63(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(30)(MULT_SIZE-1) & MULT_64(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(31)<=signed(MULT_63(31)(MULT_SIZE-1) & MULT_63(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(31)(MULT_SIZE-1) & MULT_64(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(32)<=signed(MULT_63(32)(MULT_SIZE-1) & MULT_63(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(32)(MULT_SIZE-1) & MULT_64(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(33)<=signed(MULT_63(33)(MULT_SIZE-1) & MULT_63(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(33)(MULT_SIZE-1) & MULT_64(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(34)<=signed(MULT_63(34)(MULT_SIZE-1) & MULT_63(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(34)(MULT_SIZE-1) & MULT_64(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(35)<=signed(MULT_63(35)(MULT_SIZE-1) & MULT_63(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(35)(MULT_SIZE-1) & MULT_64(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(36)<=signed(MULT_63(36)(MULT_SIZE-1) & MULT_63(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(36)(MULT_SIZE-1) & MULT_64(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(37)<=signed(MULT_63(37)(MULT_SIZE-1) & MULT_63(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(37)(MULT_SIZE-1) & MULT_64(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(38)<=signed(MULT_63(38)(MULT_SIZE-1) & MULT_63(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(38)(MULT_SIZE-1) & MULT_64(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(39)<=signed(MULT_63(39)(MULT_SIZE-1) & MULT_63(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(39)(MULT_SIZE-1) & MULT_64(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(40)<=signed(MULT_63(40)(MULT_SIZE-1) & MULT_63(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(40)(MULT_SIZE-1) & MULT_64(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(41)<=signed(MULT_63(41)(MULT_SIZE-1) & MULT_63(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(41)(MULT_SIZE-1) & MULT_64(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(42)<=signed(MULT_63(42)(MULT_SIZE-1) & MULT_63(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(42)(MULT_SIZE-1) & MULT_64(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(43)<=signed(MULT_63(43)(MULT_SIZE-1) & MULT_63(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(43)(MULT_SIZE-1) & MULT_64(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(44)<=signed(MULT_63(44)(MULT_SIZE-1) & MULT_63(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(44)(MULT_SIZE-1) & MULT_64(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(45)<=signed(MULT_63(45)(MULT_SIZE-1) & MULT_63(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(45)(MULT_SIZE-1) & MULT_64(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(46)<=signed(MULT_63(46)(MULT_SIZE-1) & MULT_63(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(46)(MULT_SIZE-1) & MULT_64(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(47)<=signed(MULT_63(47)(MULT_SIZE-1) & MULT_63(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(47)(MULT_SIZE-1) & MULT_64(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(48)<=signed(MULT_63(48)(MULT_SIZE-1) & MULT_63(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(48)(MULT_SIZE-1) & MULT_64(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(49)<=signed(MULT_63(49)(MULT_SIZE-1) & MULT_63(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(49)(MULT_SIZE-1) & MULT_64(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(50)<=signed(MULT_63(50)(MULT_SIZE-1) & MULT_63(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(50)(MULT_SIZE-1) & MULT_64(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(51)<=signed(MULT_63(51)(MULT_SIZE-1) & MULT_63(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(51)(MULT_SIZE-1) & MULT_64(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(52)<=signed(MULT_63(52)(MULT_SIZE-1) & MULT_63(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(52)(MULT_SIZE-1) & MULT_64(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(53)<=signed(MULT_63(53)(MULT_SIZE-1) & MULT_63(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(53)(MULT_SIZE-1) & MULT_64(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(54)<=signed(MULT_63(54)(MULT_SIZE-1) & MULT_63(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(54)(MULT_SIZE-1) & MULT_64(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(55)<=signed(MULT_63(55)(MULT_SIZE-1) & MULT_63(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(55)(MULT_SIZE-1) & MULT_64(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(56)<=signed(MULT_63(56)(MULT_SIZE-1) & MULT_63(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(56)(MULT_SIZE-1) & MULT_64(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(57)<=signed(MULT_63(57)(MULT_SIZE-1) & MULT_63(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(57)(MULT_SIZE-1) & MULT_64(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(58)<=signed(MULT_63(58)(MULT_SIZE-1) & MULT_63(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(58)(MULT_SIZE-1) & MULT_64(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(59)<=signed(MULT_63(59)(MULT_SIZE-1) & MULT_63(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(59)(MULT_SIZE-1) & MULT_64(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(60)<=signed(MULT_63(60)(MULT_SIZE-1) & MULT_63(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(60)(MULT_SIZE-1) & MULT_64(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(61)<=signed(MULT_63(61)(MULT_SIZE-1) & MULT_63(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(61)(MULT_SIZE-1) & MULT_64(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(62)<=signed(MULT_63(62)(MULT_SIZE-1) & MULT_63(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(62)(MULT_SIZE-1) & MULT_64(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(63)<=signed(MULT_63(63)(MULT_SIZE-1) & MULT_63(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(63)(MULT_SIZE-1) & MULT_64(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(64)<=signed(MULT_63(64)(MULT_SIZE-1) & MULT_63(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(64)(MULT_SIZE-1) & MULT_64(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(65)<=signed(MULT_63(65)(MULT_SIZE-1) & MULT_63(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(65)(MULT_SIZE-1) & MULT_64(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(66)<=signed(MULT_63(66)(MULT_SIZE-1) & MULT_63(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(66)(MULT_SIZE-1) & MULT_64(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(67)<=signed(MULT_63(67)(MULT_SIZE-1) & MULT_63(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(67)(MULT_SIZE-1) & MULT_64(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(68)<=signed(MULT_63(68)(MULT_SIZE-1) & MULT_63(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(68)(MULT_SIZE-1) & MULT_64(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(69)<=signed(MULT_63(69)(MULT_SIZE-1) & MULT_63(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(69)(MULT_SIZE-1) & MULT_64(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(70)<=signed(MULT_63(70)(MULT_SIZE-1) & MULT_63(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(70)(MULT_SIZE-1) & MULT_64(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(71)<=signed(MULT_63(71)(MULT_SIZE-1) & MULT_63(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(71)(MULT_SIZE-1) & MULT_64(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(72)<=signed(MULT_63(72)(MULT_SIZE-1) & MULT_63(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(72)(MULT_SIZE-1) & MULT_64(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(73)<=signed(MULT_63(73)(MULT_SIZE-1) & MULT_63(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(73)(MULT_SIZE-1) & MULT_64(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(74)<=signed(MULT_63(74)(MULT_SIZE-1) & MULT_63(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(74)(MULT_SIZE-1) & MULT_64(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(75)<=signed(MULT_63(75)(MULT_SIZE-1) & MULT_63(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(75)(MULT_SIZE-1) & MULT_64(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(76)<=signed(MULT_63(76)(MULT_SIZE-1) & MULT_63(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(76)(MULT_SIZE-1) & MULT_64(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(77)<=signed(MULT_63(77)(MULT_SIZE-1) & MULT_63(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(77)(MULT_SIZE-1) & MULT_64(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(78)<=signed(MULT_63(78)(MULT_SIZE-1) & MULT_63(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(78)(MULT_SIZE-1) & MULT_64(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(79)<=signed(MULT_63(79)(MULT_SIZE-1) & MULT_63(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(79)(MULT_SIZE-1) & MULT_64(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(80)<=signed(MULT_63(80)(MULT_SIZE-1) & MULT_63(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(80)(MULT_SIZE-1) & MULT_64(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(81)<=signed(MULT_63(81)(MULT_SIZE-1) & MULT_63(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(81)(MULT_SIZE-1) & MULT_64(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(82)<=signed(MULT_63(82)(MULT_SIZE-1) & MULT_63(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(82)(MULT_SIZE-1) & MULT_64(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_32(83)<=signed(MULT_63(83)(MULT_SIZE-1) & MULT_63(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_64(83)(MULT_SIZE-1) & MULT_64(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_33(0)<=signed(MULT_65(0)(MULT_SIZE-1) & MULT_65(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(0)(MULT_SIZE-1) & MULT_66(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(1)<=signed(MULT_65(1)(MULT_SIZE-1) & MULT_65(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(1)(MULT_SIZE-1) & MULT_66(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(2)<=signed(MULT_65(2)(MULT_SIZE-1) & MULT_65(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(2)(MULT_SIZE-1) & MULT_66(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(3)<=signed(MULT_65(3)(MULT_SIZE-1) & MULT_65(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(3)(MULT_SIZE-1) & MULT_66(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(4)<=signed(MULT_65(4)(MULT_SIZE-1) & MULT_65(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(4)(MULT_SIZE-1) & MULT_66(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(5)<=signed(MULT_65(5)(MULT_SIZE-1) & MULT_65(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(5)(MULT_SIZE-1) & MULT_66(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(6)<=signed(MULT_65(6)(MULT_SIZE-1) & MULT_65(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(6)(MULT_SIZE-1) & MULT_66(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(7)<=signed(MULT_65(7)(MULT_SIZE-1) & MULT_65(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(7)(MULT_SIZE-1) & MULT_66(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(8)<=signed(MULT_65(8)(MULT_SIZE-1) & MULT_65(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(8)(MULT_SIZE-1) & MULT_66(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(9)<=signed(MULT_65(9)(MULT_SIZE-1) & MULT_65(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(9)(MULT_SIZE-1) & MULT_66(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(10)<=signed(MULT_65(10)(MULT_SIZE-1) & MULT_65(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(10)(MULT_SIZE-1) & MULT_66(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(11)<=signed(MULT_65(11)(MULT_SIZE-1) & MULT_65(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(11)(MULT_SIZE-1) & MULT_66(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(12)<=signed(MULT_65(12)(MULT_SIZE-1) & MULT_65(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(12)(MULT_SIZE-1) & MULT_66(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(13)<=signed(MULT_65(13)(MULT_SIZE-1) & MULT_65(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(13)(MULT_SIZE-1) & MULT_66(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(14)<=signed(MULT_65(14)(MULT_SIZE-1) & MULT_65(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(14)(MULT_SIZE-1) & MULT_66(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(15)<=signed(MULT_65(15)(MULT_SIZE-1) & MULT_65(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(15)(MULT_SIZE-1) & MULT_66(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(16)<=signed(MULT_65(16)(MULT_SIZE-1) & MULT_65(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(16)(MULT_SIZE-1) & MULT_66(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(17)<=signed(MULT_65(17)(MULT_SIZE-1) & MULT_65(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(17)(MULT_SIZE-1) & MULT_66(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(18)<=signed(MULT_65(18)(MULT_SIZE-1) & MULT_65(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(18)(MULT_SIZE-1) & MULT_66(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(19)<=signed(MULT_65(19)(MULT_SIZE-1) & MULT_65(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(19)(MULT_SIZE-1) & MULT_66(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(20)<=signed(MULT_65(20)(MULT_SIZE-1) & MULT_65(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(20)(MULT_SIZE-1) & MULT_66(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(21)<=signed(MULT_65(21)(MULT_SIZE-1) & MULT_65(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(21)(MULT_SIZE-1) & MULT_66(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(22)<=signed(MULT_65(22)(MULT_SIZE-1) & MULT_65(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(22)(MULT_SIZE-1) & MULT_66(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(23)<=signed(MULT_65(23)(MULT_SIZE-1) & MULT_65(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(23)(MULT_SIZE-1) & MULT_66(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(24)<=signed(MULT_65(24)(MULT_SIZE-1) & MULT_65(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(24)(MULT_SIZE-1) & MULT_66(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(25)<=signed(MULT_65(25)(MULT_SIZE-1) & MULT_65(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(25)(MULT_SIZE-1) & MULT_66(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(26)<=signed(MULT_65(26)(MULT_SIZE-1) & MULT_65(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(26)(MULT_SIZE-1) & MULT_66(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(27)<=signed(MULT_65(27)(MULT_SIZE-1) & MULT_65(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(27)(MULT_SIZE-1) & MULT_66(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(28)<=signed(MULT_65(28)(MULT_SIZE-1) & MULT_65(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(28)(MULT_SIZE-1) & MULT_66(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(29)<=signed(MULT_65(29)(MULT_SIZE-1) & MULT_65(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(29)(MULT_SIZE-1) & MULT_66(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(30)<=signed(MULT_65(30)(MULT_SIZE-1) & MULT_65(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(30)(MULT_SIZE-1) & MULT_66(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(31)<=signed(MULT_65(31)(MULT_SIZE-1) & MULT_65(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(31)(MULT_SIZE-1) & MULT_66(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(32)<=signed(MULT_65(32)(MULT_SIZE-1) & MULT_65(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(32)(MULT_SIZE-1) & MULT_66(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(33)<=signed(MULT_65(33)(MULT_SIZE-1) & MULT_65(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(33)(MULT_SIZE-1) & MULT_66(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(34)<=signed(MULT_65(34)(MULT_SIZE-1) & MULT_65(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(34)(MULT_SIZE-1) & MULT_66(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(35)<=signed(MULT_65(35)(MULT_SIZE-1) & MULT_65(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(35)(MULT_SIZE-1) & MULT_66(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(36)<=signed(MULT_65(36)(MULT_SIZE-1) & MULT_65(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(36)(MULT_SIZE-1) & MULT_66(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(37)<=signed(MULT_65(37)(MULT_SIZE-1) & MULT_65(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(37)(MULT_SIZE-1) & MULT_66(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(38)<=signed(MULT_65(38)(MULT_SIZE-1) & MULT_65(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(38)(MULT_SIZE-1) & MULT_66(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(39)<=signed(MULT_65(39)(MULT_SIZE-1) & MULT_65(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(39)(MULT_SIZE-1) & MULT_66(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(40)<=signed(MULT_65(40)(MULT_SIZE-1) & MULT_65(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(40)(MULT_SIZE-1) & MULT_66(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(41)<=signed(MULT_65(41)(MULT_SIZE-1) & MULT_65(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(41)(MULT_SIZE-1) & MULT_66(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(42)<=signed(MULT_65(42)(MULT_SIZE-1) & MULT_65(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(42)(MULT_SIZE-1) & MULT_66(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(43)<=signed(MULT_65(43)(MULT_SIZE-1) & MULT_65(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(43)(MULT_SIZE-1) & MULT_66(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(44)<=signed(MULT_65(44)(MULT_SIZE-1) & MULT_65(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(44)(MULT_SIZE-1) & MULT_66(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(45)<=signed(MULT_65(45)(MULT_SIZE-1) & MULT_65(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(45)(MULT_SIZE-1) & MULT_66(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(46)<=signed(MULT_65(46)(MULT_SIZE-1) & MULT_65(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(46)(MULT_SIZE-1) & MULT_66(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(47)<=signed(MULT_65(47)(MULT_SIZE-1) & MULT_65(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(47)(MULT_SIZE-1) & MULT_66(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(48)<=signed(MULT_65(48)(MULT_SIZE-1) & MULT_65(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(48)(MULT_SIZE-1) & MULT_66(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(49)<=signed(MULT_65(49)(MULT_SIZE-1) & MULT_65(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(49)(MULT_SIZE-1) & MULT_66(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(50)<=signed(MULT_65(50)(MULT_SIZE-1) & MULT_65(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(50)(MULT_SIZE-1) & MULT_66(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(51)<=signed(MULT_65(51)(MULT_SIZE-1) & MULT_65(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(51)(MULT_SIZE-1) & MULT_66(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(52)<=signed(MULT_65(52)(MULT_SIZE-1) & MULT_65(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(52)(MULT_SIZE-1) & MULT_66(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(53)<=signed(MULT_65(53)(MULT_SIZE-1) & MULT_65(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(53)(MULT_SIZE-1) & MULT_66(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(54)<=signed(MULT_65(54)(MULT_SIZE-1) & MULT_65(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(54)(MULT_SIZE-1) & MULT_66(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(55)<=signed(MULT_65(55)(MULT_SIZE-1) & MULT_65(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(55)(MULT_SIZE-1) & MULT_66(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(56)<=signed(MULT_65(56)(MULT_SIZE-1) & MULT_65(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(56)(MULT_SIZE-1) & MULT_66(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(57)<=signed(MULT_65(57)(MULT_SIZE-1) & MULT_65(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(57)(MULT_SIZE-1) & MULT_66(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(58)<=signed(MULT_65(58)(MULT_SIZE-1) & MULT_65(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(58)(MULT_SIZE-1) & MULT_66(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(59)<=signed(MULT_65(59)(MULT_SIZE-1) & MULT_65(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(59)(MULT_SIZE-1) & MULT_66(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(60)<=signed(MULT_65(60)(MULT_SIZE-1) & MULT_65(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(60)(MULT_SIZE-1) & MULT_66(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(61)<=signed(MULT_65(61)(MULT_SIZE-1) & MULT_65(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(61)(MULT_SIZE-1) & MULT_66(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(62)<=signed(MULT_65(62)(MULT_SIZE-1) & MULT_65(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(62)(MULT_SIZE-1) & MULT_66(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(63)<=signed(MULT_65(63)(MULT_SIZE-1) & MULT_65(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(63)(MULT_SIZE-1) & MULT_66(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(64)<=signed(MULT_65(64)(MULT_SIZE-1) & MULT_65(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(64)(MULT_SIZE-1) & MULT_66(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(65)<=signed(MULT_65(65)(MULT_SIZE-1) & MULT_65(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(65)(MULT_SIZE-1) & MULT_66(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(66)<=signed(MULT_65(66)(MULT_SIZE-1) & MULT_65(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(66)(MULT_SIZE-1) & MULT_66(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(67)<=signed(MULT_65(67)(MULT_SIZE-1) & MULT_65(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(67)(MULT_SIZE-1) & MULT_66(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(68)<=signed(MULT_65(68)(MULT_SIZE-1) & MULT_65(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(68)(MULT_SIZE-1) & MULT_66(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(69)<=signed(MULT_65(69)(MULT_SIZE-1) & MULT_65(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(69)(MULT_SIZE-1) & MULT_66(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(70)<=signed(MULT_65(70)(MULT_SIZE-1) & MULT_65(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(70)(MULT_SIZE-1) & MULT_66(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(71)<=signed(MULT_65(71)(MULT_SIZE-1) & MULT_65(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(71)(MULT_SIZE-1) & MULT_66(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(72)<=signed(MULT_65(72)(MULT_SIZE-1) & MULT_65(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(72)(MULT_SIZE-1) & MULT_66(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(73)<=signed(MULT_65(73)(MULT_SIZE-1) & MULT_65(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(73)(MULT_SIZE-1) & MULT_66(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(74)<=signed(MULT_65(74)(MULT_SIZE-1) & MULT_65(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(74)(MULT_SIZE-1) & MULT_66(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(75)<=signed(MULT_65(75)(MULT_SIZE-1) & MULT_65(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(75)(MULT_SIZE-1) & MULT_66(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(76)<=signed(MULT_65(76)(MULT_SIZE-1) & MULT_65(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(76)(MULT_SIZE-1) & MULT_66(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(77)<=signed(MULT_65(77)(MULT_SIZE-1) & MULT_65(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(77)(MULT_SIZE-1) & MULT_66(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(78)<=signed(MULT_65(78)(MULT_SIZE-1) & MULT_65(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(78)(MULT_SIZE-1) & MULT_66(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(79)<=signed(MULT_65(79)(MULT_SIZE-1) & MULT_65(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(79)(MULT_SIZE-1) & MULT_66(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(80)<=signed(MULT_65(80)(MULT_SIZE-1) & MULT_65(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(80)(MULT_SIZE-1) & MULT_66(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(81)<=signed(MULT_65(81)(MULT_SIZE-1) & MULT_65(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(81)(MULT_SIZE-1) & MULT_66(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(82)<=signed(MULT_65(82)(MULT_SIZE-1) & MULT_65(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(82)(MULT_SIZE-1) & MULT_66(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_33(83)<=signed(MULT_65(83)(MULT_SIZE-1) & MULT_65(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_66(83)(MULT_SIZE-1) & MULT_66(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_34(0)<=signed(MULT_67(0)(MULT_SIZE-1) & MULT_67(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(0)(MULT_SIZE-1) & MULT_68(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(1)<=signed(MULT_67(1)(MULT_SIZE-1) & MULT_67(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(1)(MULT_SIZE-1) & MULT_68(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(2)<=signed(MULT_67(2)(MULT_SIZE-1) & MULT_67(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(2)(MULT_SIZE-1) & MULT_68(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(3)<=signed(MULT_67(3)(MULT_SIZE-1) & MULT_67(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(3)(MULT_SIZE-1) & MULT_68(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(4)<=signed(MULT_67(4)(MULT_SIZE-1) & MULT_67(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(4)(MULT_SIZE-1) & MULT_68(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(5)<=signed(MULT_67(5)(MULT_SIZE-1) & MULT_67(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(5)(MULT_SIZE-1) & MULT_68(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(6)<=signed(MULT_67(6)(MULT_SIZE-1) & MULT_67(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(6)(MULT_SIZE-1) & MULT_68(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(7)<=signed(MULT_67(7)(MULT_SIZE-1) & MULT_67(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(7)(MULT_SIZE-1) & MULT_68(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(8)<=signed(MULT_67(8)(MULT_SIZE-1) & MULT_67(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(8)(MULT_SIZE-1) & MULT_68(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(9)<=signed(MULT_67(9)(MULT_SIZE-1) & MULT_67(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(9)(MULT_SIZE-1) & MULT_68(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(10)<=signed(MULT_67(10)(MULT_SIZE-1) & MULT_67(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(10)(MULT_SIZE-1) & MULT_68(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(11)<=signed(MULT_67(11)(MULT_SIZE-1) & MULT_67(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(11)(MULT_SIZE-1) & MULT_68(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(12)<=signed(MULT_67(12)(MULT_SIZE-1) & MULT_67(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(12)(MULT_SIZE-1) & MULT_68(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(13)<=signed(MULT_67(13)(MULT_SIZE-1) & MULT_67(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(13)(MULT_SIZE-1) & MULT_68(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(14)<=signed(MULT_67(14)(MULT_SIZE-1) & MULT_67(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(14)(MULT_SIZE-1) & MULT_68(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(15)<=signed(MULT_67(15)(MULT_SIZE-1) & MULT_67(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(15)(MULT_SIZE-1) & MULT_68(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(16)<=signed(MULT_67(16)(MULT_SIZE-1) & MULT_67(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(16)(MULT_SIZE-1) & MULT_68(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(17)<=signed(MULT_67(17)(MULT_SIZE-1) & MULT_67(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(17)(MULT_SIZE-1) & MULT_68(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(18)<=signed(MULT_67(18)(MULT_SIZE-1) & MULT_67(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(18)(MULT_SIZE-1) & MULT_68(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(19)<=signed(MULT_67(19)(MULT_SIZE-1) & MULT_67(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(19)(MULT_SIZE-1) & MULT_68(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(20)<=signed(MULT_67(20)(MULT_SIZE-1) & MULT_67(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(20)(MULT_SIZE-1) & MULT_68(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(21)<=signed(MULT_67(21)(MULT_SIZE-1) & MULT_67(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(21)(MULT_SIZE-1) & MULT_68(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(22)<=signed(MULT_67(22)(MULT_SIZE-1) & MULT_67(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(22)(MULT_SIZE-1) & MULT_68(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(23)<=signed(MULT_67(23)(MULT_SIZE-1) & MULT_67(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(23)(MULT_SIZE-1) & MULT_68(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(24)<=signed(MULT_67(24)(MULT_SIZE-1) & MULT_67(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(24)(MULT_SIZE-1) & MULT_68(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(25)<=signed(MULT_67(25)(MULT_SIZE-1) & MULT_67(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(25)(MULT_SIZE-1) & MULT_68(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(26)<=signed(MULT_67(26)(MULT_SIZE-1) & MULT_67(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(26)(MULT_SIZE-1) & MULT_68(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(27)<=signed(MULT_67(27)(MULT_SIZE-1) & MULT_67(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(27)(MULT_SIZE-1) & MULT_68(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(28)<=signed(MULT_67(28)(MULT_SIZE-1) & MULT_67(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(28)(MULT_SIZE-1) & MULT_68(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(29)<=signed(MULT_67(29)(MULT_SIZE-1) & MULT_67(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(29)(MULT_SIZE-1) & MULT_68(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(30)<=signed(MULT_67(30)(MULT_SIZE-1) & MULT_67(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(30)(MULT_SIZE-1) & MULT_68(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(31)<=signed(MULT_67(31)(MULT_SIZE-1) & MULT_67(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(31)(MULT_SIZE-1) & MULT_68(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(32)<=signed(MULT_67(32)(MULT_SIZE-1) & MULT_67(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(32)(MULT_SIZE-1) & MULT_68(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(33)<=signed(MULT_67(33)(MULT_SIZE-1) & MULT_67(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(33)(MULT_SIZE-1) & MULT_68(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(34)<=signed(MULT_67(34)(MULT_SIZE-1) & MULT_67(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(34)(MULT_SIZE-1) & MULT_68(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(35)<=signed(MULT_67(35)(MULT_SIZE-1) & MULT_67(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(35)(MULT_SIZE-1) & MULT_68(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(36)<=signed(MULT_67(36)(MULT_SIZE-1) & MULT_67(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(36)(MULT_SIZE-1) & MULT_68(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(37)<=signed(MULT_67(37)(MULT_SIZE-1) & MULT_67(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(37)(MULT_SIZE-1) & MULT_68(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(38)<=signed(MULT_67(38)(MULT_SIZE-1) & MULT_67(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(38)(MULT_SIZE-1) & MULT_68(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(39)<=signed(MULT_67(39)(MULT_SIZE-1) & MULT_67(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(39)(MULT_SIZE-1) & MULT_68(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(40)<=signed(MULT_67(40)(MULT_SIZE-1) & MULT_67(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(40)(MULT_SIZE-1) & MULT_68(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(41)<=signed(MULT_67(41)(MULT_SIZE-1) & MULT_67(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(41)(MULT_SIZE-1) & MULT_68(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(42)<=signed(MULT_67(42)(MULT_SIZE-1) & MULT_67(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(42)(MULT_SIZE-1) & MULT_68(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(43)<=signed(MULT_67(43)(MULT_SIZE-1) & MULT_67(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(43)(MULT_SIZE-1) & MULT_68(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(44)<=signed(MULT_67(44)(MULT_SIZE-1) & MULT_67(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(44)(MULT_SIZE-1) & MULT_68(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(45)<=signed(MULT_67(45)(MULT_SIZE-1) & MULT_67(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(45)(MULT_SIZE-1) & MULT_68(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(46)<=signed(MULT_67(46)(MULT_SIZE-1) & MULT_67(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(46)(MULT_SIZE-1) & MULT_68(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(47)<=signed(MULT_67(47)(MULT_SIZE-1) & MULT_67(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(47)(MULT_SIZE-1) & MULT_68(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(48)<=signed(MULT_67(48)(MULT_SIZE-1) & MULT_67(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(48)(MULT_SIZE-1) & MULT_68(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(49)<=signed(MULT_67(49)(MULT_SIZE-1) & MULT_67(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(49)(MULT_SIZE-1) & MULT_68(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(50)<=signed(MULT_67(50)(MULT_SIZE-1) & MULT_67(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(50)(MULT_SIZE-1) & MULT_68(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(51)<=signed(MULT_67(51)(MULT_SIZE-1) & MULT_67(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(51)(MULT_SIZE-1) & MULT_68(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(52)<=signed(MULT_67(52)(MULT_SIZE-1) & MULT_67(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(52)(MULT_SIZE-1) & MULT_68(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(53)<=signed(MULT_67(53)(MULT_SIZE-1) & MULT_67(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(53)(MULT_SIZE-1) & MULT_68(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(54)<=signed(MULT_67(54)(MULT_SIZE-1) & MULT_67(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(54)(MULT_SIZE-1) & MULT_68(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(55)<=signed(MULT_67(55)(MULT_SIZE-1) & MULT_67(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(55)(MULT_SIZE-1) & MULT_68(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(56)<=signed(MULT_67(56)(MULT_SIZE-1) & MULT_67(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(56)(MULT_SIZE-1) & MULT_68(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(57)<=signed(MULT_67(57)(MULT_SIZE-1) & MULT_67(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(57)(MULT_SIZE-1) & MULT_68(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(58)<=signed(MULT_67(58)(MULT_SIZE-1) & MULT_67(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(58)(MULT_SIZE-1) & MULT_68(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(59)<=signed(MULT_67(59)(MULT_SIZE-1) & MULT_67(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(59)(MULT_SIZE-1) & MULT_68(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(60)<=signed(MULT_67(60)(MULT_SIZE-1) & MULT_67(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(60)(MULT_SIZE-1) & MULT_68(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(61)<=signed(MULT_67(61)(MULT_SIZE-1) & MULT_67(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(61)(MULT_SIZE-1) & MULT_68(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(62)<=signed(MULT_67(62)(MULT_SIZE-1) & MULT_67(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(62)(MULT_SIZE-1) & MULT_68(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(63)<=signed(MULT_67(63)(MULT_SIZE-1) & MULT_67(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(63)(MULT_SIZE-1) & MULT_68(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(64)<=signed(MULT_67(64)(MULT_SIZE-1) & MULT_67(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(64)(MULT_SIZE-1) & MULT_68(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(65)<=signed(MULT_67(65)(MULT_SIZE-1) & MULT_67(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(65)(MULT_SIZE-1) & MULT_68(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(66)<=signed(MULT_67(66)(MULT_SIZE-1) & MULT_67(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(66)(MULT_SIZE-1) & MULT_68(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(67)<=signed(MULT_67(67)(MULT_SIZE-1) & MULT_67(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(67)(MULT_SIZE-1) & MULT_68(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(68)<=signed(MULT_67(68)(MULT_SIZE-1) & MULT_67(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(68)(MULT_SIZE-1) & MULT_68(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(69)<=signed(MULT_67(69)(MULT_SIZE-1) & MULT_67(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(69)(MULT_SIZE-1) & MULT_68(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(70)<=signed(MULT_67(70)(MULT_SIZE-1) & MULT_67(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(70)(MULT_SIZE-1) & MULT_68(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(71)<=signed(MULT_67(71)(MULT_SIZE-1) & MULT_67(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(71)(MULT_SIZE-1) & MULT_68(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(72)<=signed(MULT_67(72)(MULT_SIZE-1) & MULT_67(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(72)(MULT_SIZE-1) & MULT_68(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(73)<=signed(MULT_67(73)(MULT_SIZE-1) & MULT_67(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(73)(MULT_SIZE-1) & MULT_68(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(74)<=signed(MULT_67(74)(MULT_SIZE-1) & MULT_67(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(74)(MULT_SIZE-1) & MULT_68(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(75)<=signed(MULT_67(75)(MULT_SIZE-1) & MULT_67(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(75)(MULT_SIZE-1) & MULT_68(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(76)<=signed(MULT_67(76)(MULT_SIZE-1) & MULT_67(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(76)(MULT_SIZE-1) & MULT_68(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(77)<=signed(MULT_67(77)(MULT_SIZE-1) & MULT_67(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(77)(MULT_SIZE-1) & MULT_68(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(78)<=signed(MULT_67(78)(MULT_SIZE-1) & MULT_67(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(78)(MULT_SIZE-1) & MULT_68(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(79)<=signed(MULT_67(79)(MULT_SIZE-1) & MULT_67(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(79)(MULT_SIZE-1) & MULT_68(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(80)<=signed(MULT_67(80)(MULT_SIZE-1) & MULT_67(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(80)(MULT_SIZE-1) & MULT_68(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(81)<=signed(MULT_67(81)(MULT_SIZE-1) & MULT_67(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(81)(MULT_SIZE-1) & MULT_68(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(82)<=signed(MULT_67(82)(MULT_SIZE-1) & MULT_67(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(82)(MULT_SIZE-1) & MULT_68(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_34(83)<=signed(MULT_67(83)(MULT_SIZE-1) & MULT_67(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_68(83)(MULT_SIZE-1) & MULT_68(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_35(0)<=signed(MULT_69(0)(MULT_SIZE-1) & MULT_69(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(0)(MULT_SIZE-1) & MULT_70(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(1)<=signed(MULT_69(1)(MULT_SIZE-1) & MULT_69(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(1)(MULT_SIZE-1) & MULT_70(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(2)<=signed(MULT_69(2)(MULT_SIZE-1) & MULT_69(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(2)(MULT_SIZE-1) & MULT_70(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(3)<=signed(MULT_69(3)(MULT_SIZE-1) & MULT_69(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(3)(MULT_SIZE-1) & MULT_70(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(4)<=signed(MULT_69(4)(MULT_SIZE-1) & MULT_69(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(4)(MULT_SIZE-1) & MULT_70(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(5)<=signed(MULT_69(5)(MULT_SIZE-1) & MULT_69(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(5)(MULT_SIZE-1) & MULT_70(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(6)<=signed(MULT_69(6)(MULT_SIZE-1) & MULT_69(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(6)(MULT_SIZE-1) & MULT_70(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(7)<=signed(MULT_69(7)(MULT_SIZE-1) & MULT_69(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(7)(MULT_SIZE-1) & MULT_70(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(8)<=signed(MULT_69(8)(MULT_SIZE-1) & MULT_69(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(8)(MULT_SIZE-1) & MULT_70(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(9)<=signed(MULT_69(9)(MULT_SIZE-1) & MULT_69(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(9)(MULT_SIZE-1) & MULT_70(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(10)<=signed(MULT_69(10)(MULT_SIZE-1) & MULT_69(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(10)(MULT_SIZE-1) & MULT_70(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(11)<=signed(MULT_69(11)(MULT_SIZE-1) & MULT_69(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(11)(MULT_SIZE-1) & MULT_70(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(12)<=signed(MULT_69(12)(MULT_SIZE-1) & MULT_69(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(12)(MULT_SIZE-1) & MULT_70(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(13)<=signed(MULT_69(13)(MULT_SIZE-1) & MULT_69(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(13)(MULT_SIZE-1) & MULT_70(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(14)<=signed(MULT_69(14)(MULT_SIZE-1) & MULT_69(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(14)(MULT_SIZE-1) & MULT_70(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(15)<=signed(MULT_69(15)(MULT_SIZE-1) & MULT_69(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(15)(MULT_SIZE-1) & MULT_70(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(16)<=signed(MULT_69(16)(MULT_SIZE-1) & MULT_69(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(16)(MULT_SIZE-1) & MULT_70(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(17)<=signed(MULT_69(17)(MULT_SIZE-1) & MULT_69(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(17)(MULT_SIZE-1) & MULT_70(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(18)<=signed(MULT_69(18)(MULT_SIZE-1) & MULT_69(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(18)(MULT_SIZE-1) & MULT_70(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(19)<=signed(MULT_69(19)(MULT_SIZE-1) & MULT_69(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(19)(MULT_SIZE-1) & MULT_70(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(20)<=signed(MULT_69(20)(MULT_SIZE-1) & MULT_69(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(20)(MULT_SIZE-1) & MULT_70(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(21)<=signed(MULT_69(21)(MULT_SIZE-1) & MULT_69(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(21)(MULT_SIZE-1) & MULT_70(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(22)<=signed(MULT_69(22)(MULT_SIZE-1) & MULT_69(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(22)(MULT_SIZE-1) & MULT_70(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(23)<=signed(MULT_69(23)(MULT_SIZE-1) & MULT_69(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(23)(MULT_SIZE-1) & MULT_70(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(24)<=signed(MULT_69(24)(MULT_SIZE-1) & MULT_69(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(24)(MULT_SIZE-1) & MULT_70(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(25)<=signed(MULT_69(25)(MULT_SIZE-1) & MULT_69(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(25)(MULT_SIZE-1) & MULT_70(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(26)<=signed(MULT_69(26)(MULT_SIZE-1) & MULT_69(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(26)(MULT_SIZE-1) & MULT_70(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(27)<=signed(MULT_69(27)(MULT_SIZE-1) & MULT_69(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(27)(MULT_SIZE-1) & MULT_70(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(28)<=signed(MULT_69(28)(MULT_SIZE-1) & MULT_69(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(28)(MULT_SIZE-1) & MULT_70(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(29)<=signed(MULT_69(29)(MULT_SIZE-1) & MULT_69(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(29)(MULT_SIZE-1) & MULT_70(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(30)<=signed(MULT_69(30)(MULT_SIZE-1) & MULT_69(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(30)(MULT_SIZE-1) & MULT_70(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(31)<=signed(MULT_69(31)(MULT_SIZE-1) & MULT_69(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(31)(MULT_SIZE-1) & MULT_70(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(32)<=signed(MULT_69(32)(MULT_SIZE-1) & MULT_69(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(32)(MULT_SIZE-1) & MULT_70(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(33)<=signed(MULT_69(33)(MULT_SIZE-1) & MULT_69(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(33)(MULT_SIZE-1) & MULT_70(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(34)<=signed(MULT_69(34)(MULT_SIZE-1) & MULT_69(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(34)(MULT_SIZE-1) & MULT_70(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(35)<=signed(MULT_69(35)(MULT_SIZE-1) & MULT_69(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(35)(MULT_SIZE-1) & MULT_70(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(36)<=signed(MULT_69(36)(MULT_SIZE-1) & MULT_69(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(36)(MULT_SIZE-1) & MULT_70(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(37)<=signed(MULT_69(37)(MULT_SIZE-1) & MULT_69(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(37)(MULT_SIZE-1) & MULT_70(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(38)<=signed(MULT_69(38)(MULT_SIZE-1) & MULT_69(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(38)(MULT_SIZE-1) & MULT_70(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(39)<=signed(MULT_69(39)(MULT_SIZE-1) & MULT_69(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(39)(MULT_SIZE-1) & MULT_70(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(40)<=signed(MULT_69(40)(MULT_SIZE-1) & MULT_69(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(40)(MULT_SIZE-1) & MULT_70(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(41)<=signed(MULT_69(41)(MULT_SIZE-1) & MULT_69(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(41)(MULT_SIZE-1) & MULT_70(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(42)<=signed(MULT_69(42)(MULT_SIZE-1) & MULT_69(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(42)(MULT_SIZE-1) & MULT_70(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(43)<=signed(MULT_69(43)(MULT_SIZE-1) & MULT_69(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(43)(MULT_SIZE-1) & MULT_70(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(44)<=signed(MULT_69(44)(MULT_SIZE-1) & MULT_69(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(44)(MULT_SIZE-1) & MULT_70(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(45)<=signed(MULT_69(45)(MULT_SIZE-1) & MULT_69(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(45)(MULT_SIZE-1) & MULT_70(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(46)<=signed(MULT_69(46)(MULT_SIZE-1) & MULT_69(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(46)(MULT_SIZE-1) & MULT_70(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(47)<=signed(MULT_69(47)(MULT_SIZE-1) & MULT_69(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(47)(MULT_SIZE-1) & MULT_70(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(48)<=signed(MULT_69(48)(MULT_SIZE-1) & MULT_69(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(48)(MULT_SIZE-1) & MULT_70(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(49)<=signed(MULT_69(49)(MULT_SIZE-1) & MULT_69(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(49)(MULT_SIZE-1) & MULT_70(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(50)<=signed(MULT_69(50)(MULT_SIZE-1) & MULT_69(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(50)(MULT_SIZE-1) & MULT_70(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(51)<=signed(MULT_69(51)(MULT_SIZE-1) & MULT_69(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(51)(MULT_SIZE-1) & MULT_70(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(52)<=signed(MULT_69(52)(MULT_SIZE-1) & MULT_69(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(52)(MULT_SIZE-1) & MULT_70(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(53)<=signed(MULT_69(53)(MULT_SIZE-1) & MULT_69(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(53)(MULT_SIZE-1) & MULT_70(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(54)<=signed(MULT_69(54)(MULT_SIZE-1) & MULT_69(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(54)(MULT_SIZE-1) & MULT_70(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(55)<=signed(MULT_69(55)(MULT_SIZE-1) & MULT_69(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(55)(MULT_SIZE-1) & MULT_70(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(56)<=signed(MULT_69(56)(MULT_SIZE-1) & MULT_69(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(56)(MULT_SIZE-1) & MULT_70(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(57)<=signed(MULT_69(57)(MULT_SIZE-1) & MULT_69(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(57)(MULT_SIZE-1) & MULT_70(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(58)<=signed(MULT_69(58)(MULT_SIZE-1) & MULT_69(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(58)(MULT_SIZE-1) & MULT_70(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(59)<=signed(MULT_69(59)(MULT_SIZE-1) & MULT_69(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(59)(MULT_SIZE-1) & MULT_70(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(60)<=signed(MULT_69(60)(MULT_SIZE-1) & MULT_69(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(60)(MULT_SIZE-1) & MULT_70(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(61)<=signed(MULT_69(61)(MULT_SIZE-1) & MULT_69(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(61)(MULT_SIZE-1) & MULT_70(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(62)<=signed(MULT_69(62)(MULT_SIZE-1) & MULT_69(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(62)(MULT_SIZE-1) & MULT_70(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(63)<=signed(MULT_69(63)(MULT_SIZE-1) & MULT_69(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(63)(MULT_SIZE-1) & MULT_70(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(64)<=signed(MULT_69(64)(MULT_SIZE-1) & MULT_69(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(64)(MULT_SIZE-1) & MULT_70(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(65)<=signed(MULT_69(65)(MULT_SIZE-1) & MULT_69(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(65)(MULT_SIZE-1) & MULT_70(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(66)<=signed(MULT_69(66)(MULT_SIZE-1) & MULT_69(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(66)(MULT_SIZE-1) & MULT_70(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(67)<=signed(MULT_69(67)(MULT_SIZE-1) & MULT_69(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(67)(MULT_SIZE-1) & MULT_70(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(68)<=signed(MULT_69(68)(MULT_SIZE-1) & MULT_69(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(68)(MULT_SIZE-1) & MULT_70(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(69)<=signed(MULT_69(69)(MULT_SIZE-1) & MULT_69(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(69)(MULT_SIZE-1) & MULT_70(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(70)<=signed(MULT_69(70)(MULT_SIZE-1) & MULT_69(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(70)(MULT_SIZE-1) & MULT_70(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(71)<=signed(MULT_69(71)(MULT_SIZE-1) & MULT_69(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(71)(MULT_SIZE-1) & MULT_70(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(72)<=signed(MULT_69(72)(MULT_SIZE-1) & MULT_69(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(72)(MULT_SIZE-1) & MULT_70(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(73)<=signed(MULT_69(73)(MULT_SIZE-1) & MULT_69(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(73)(MULT_SIZE-1) & MULT_70(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(74)<=signed(MULT_69(74)(MULT_SIZE-1) & MULT_69(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(74)(MULT_SIZE-1) & MULT_70(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(75)<=signed(MULT_69(75)(MULT_SIZE-1) & MULT_69(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(75)(MULT_SIZE-1) & MULT_70(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(76)<=signed(MULT_69(76)(MULT_SIZE-1) & MULT_69(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(76)(MULT_SIZE-1) & MULT_70(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(77)<=signed(MULT_69(77)(MULT_SIZE-1) & MULT_69(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(77)(MULT_SIZE-1) & MULT_70(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(78)<=signed(MULT_69(78)(MULT_SIZE-1) & MULT_69(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(78)(MULT_SIZE-1) & MULT_70(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(79)<=signed(MULT_69(79)(MULT_SIZE-1) & MULT_69(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(79)(MULT_SIZE-1) & MULT_70(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(80)<=signed(MULT_69(80)(MULT_SIZE-1) & MULT_69(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(80)(MULT_SIZE-1) & MULT_70(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(81)<=signed(MULT_69(81)(MULT_SIZE-1) & MULT_69(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(81)(MULT_SIZE-1) & MULT_70(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(82)<=signed(MULT_69(82)(MULT_SIZE-1) & MULT_69(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(82)(MULT_SIZE-1) & MULT_70(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_35(83)<=signed(MULT_69(83)(MULT_SIZE-1) & MULT_69(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_70(83)(MULT_SIZE-1) & MULT_70(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_36(0)<=signed(MULT_71(0)(MULT_SIZE-1) & MULT_71(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(0)(MULT_SIZE-1) & MULT_72(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(1)<=signed(MULT_71(1)(MULT_SIZE-1) & MULT_71(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(1)(MULT_SIZE-1) & MULT_72(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(2)<=signed(MULT_71(2)(MULT_SIZE-1) & MULT_71(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(2)(MULT_SIZE-1) & MULT_72(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(3)<=signed(MULT_71(3)(MULT_SIZE-1) & MULT_71(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(3)(MULT_SIZE-1) & MULT_72(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(4)<=signed(MULT_71(4)(MULT_SIZE-1) & MULT_71(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(4)(MULT_SIZE-1) & MULT_72(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(5)<=signed(MULT_71(5)(MULT_SIZE-1) & MULT_71(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(5)(MULT_SIZE-1) & MULT_72(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(6)<=signed(MULT_71(6)(MULT_SIZE-1) & MULT_71(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(6)(MULT_SIZE-1) & MULT_72(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(7)<=signed(MULT_71(7)(MULT_SIZE-1) & MULT_71(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(7)(MULT_SIZE-1) & MULT_72(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(8)<=signed(MULT_71(8)(MULT_SIZE-1) & MULT_71(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(8)(MULT_SIZE-1) & MULT_72(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(9)<=signed(MULT_71(9)(MULT_SIZE-1) & MULT_71(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(9)(MULT_SIZE-1) & MULT_72(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(10)<=signed(MULT_71(10)(MULT_SIZE-1) & MULT_71(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(10)(MULT_SIZE-1) & MULT_72(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(11)<=signed(MULT_71(11)(MULT_SIZE-1) & MULT_71(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(11)(MULT_SIZE-1) & MULT_72(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(12)<=signed(MULT_71(12)(MULT_SIZE-1) & MULT_71(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(12)(MULT_SIZE-1) & MULT_72(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(13)<=signed(MULT_71(13)(MULT_SIZE-1) & MULT_71(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(13)(MULT_SIZE-1) & MULT_72(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(14)<=signed(MULT_71(14)(MULT_SIZE-1) & MULT_71(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(14)(MULT_SIZE-1) & MULT_72(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(15)<=signed(MULT_71(15)(MULT_SIZE-1) & MULT_71(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(15)(MULT_SIZE-1) & MULT_72(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(16)<=signed(MULT_71(16)(MULT_SIZE-1) & MULT_71(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(16)(MULT_SIZE-1) & MULT_72(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(17)<=signed(MULT_71(17)(MULT_SIZE-1) & MULT_71(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(17)(MULT_SIZE-1) & MULT_72(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(18)<=signed(MULT_71(18)(MULT_SIZE-1) & MULT_71(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(18)(MULT_SIZE-1) & MULT_72(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(19)<=signed(MULT_71(19)(MULT_SIZE-1) & MULT_71(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(19)(MULT_SIZE-1) & MULT_72(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(20)<=signed(MULT_71(20)(MULT_SIZE-1) & MULT_71(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(20)(MULT_SIZE-1) & MULT_72(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(21)<=signed(MULT_71(21)(MULT_SIZE-1) & MULT_71(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(21)(MULT_SIZE-1) & MULT_72(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(22)<=signed(MULT_71(22)(MULT_SIZE-1) & MULT_71(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(22)(MULT_SIZE-1) & MULT_72(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(23)<=signed(MULT_71(23)(MULT_SIZE-1) & MULT_71(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(23)(MULT_SIZE-1) & MULT_72(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(24)<=signed(MULT_71(24)(MULT_SIZE-1) & MULT_71(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(24)(MULT_SIZE-1) & MULT_72(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(25)<=signed(MULT_71(25)(MULT_SIZE-1) & MULT_71(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(25)(MULT_SIZE-1) & MULT_72(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(26)<=signed(MULT_71(26)(MULT_SIZE-1) & MULT_71(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(26)(MULT_SIZE-1) & MULT_72(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(27)<=signed(MULT_71(27)(MULT_SIZE-1) & MULT_71(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(27)(MULT_SIZE-1) & MULT_72(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(28)<=signed(MULT_71(28)(MULT_SIZE-1) & MULT_71(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(28)(MULT_SIZE-1) & MULT_72(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(29)<=signed(MULT_71(29)(MULT_SIZE-1) & MULT_71(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(29)(MULT_SIZE-1) & MULT_72(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(30)<=signed(MULT_71(30)(MULT_SIZE-1) & MULT_71(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(30)(MULT_SIZE-1) & MULT_72(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(31)<=signed(MULT_71(31)(MULT_SIZE-1) & MULT_71(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(31)(MULT_SIZE-1) & MULT_72(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(32)<=signed(MULT_71(32)(MULT_SIZE-1) & MULT_71(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(32)(MULT_SIZE-1) & MULT_72(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(33)<=signed(MULT_71(33)(MULT_SIZE-1) & MULT_71(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(33)(MULT_SIZE-1) & MULT_72(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(34)<=signed(MULT_71(34)(MULT_SIZE-1) & MULT_71(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(34)(MULT_SIZE-1) & MULT_72(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(35)<=signed(MULT_71(35)(MULT_SIZE-1) & MULT_71(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(35)(MULT_SIZE-1) & MULT_72(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(36)<=signed(MULT_71(36)(MULT_SIZE-1) & MULT_71(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(36)(MULT_SIZE-1) & MULT_72(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(37)<=signed(MULT_71(37)(MULT_SIZE-1) & MULT_71(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(37)(MULT_SIZE-1) & MULT_72(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(38)<=signed(MULT_71(38)(MULT_SIZE-1) & MULT_71(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(38)(MULT_SIZE-1) & MULT_72(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(39)<=signed(MULT_71(39)(MULT_SIZE-1) & MULT_71(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(39)(MULT_SIZE-1) & MULT_72(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(40)<=signed(MULT_71(40)(MULT_SIZE-1) & MULT_71(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(40)(MULT_SIZE-1) & MULT_72(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(41)<=signed(MULT_71(41)(MULT_SIZE-1) & MULT_71(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(41)(MULT_SIZE-1) & MULT_72(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(42)<=signed(MULT_71(42)(MULT_SIZE-1) & MULT_71(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(42)(MULT_SIZE-1) & MULT_72(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(43)<=signed(MULT_71(43)(MULT_SIZE-1) & MULT_71(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(43)(MULT_SIZE-1) & MULT_72(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(44)<=signed(MULT_71(44)(MULT_SIZE-1) & MULT_71(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(44)(MULT_SIZE-1) & MULT_72(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(45)<=signed(MULT_71(45)(MULT_SIZE-1) & MULT_71(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(45)(MULT_SIZE-1) & MULT_72(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(46)<=signed(MULT_71(46)(MULT_SIZE-1) & MULT_71(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(46)(MULT_SIZE-1) & MULT_72(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(47)<=signed(MULT_71(47)(MULT_SIZE-1) & MULT_71(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(47)(MULT_SIZE-1) & MULT_72(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(48)<=signed(MULT_71(48)(MULT_SIZE-1) & MULT_71(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(48)(MULT_SIZE-1) & MULT_72(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(49)<=signed(MULT_71(49)(MULT_SIZE-1) & MULT_71(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(49)(MULT_SIZE-1) & MULT_72(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(50)<=signed(MULT_71(50)(MULT_SIZE-1) & MULT_71(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(50)(MULT_SIZE-1) & MULT_72(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(51)<=signed(MULT_71(51)(MULT_SIZE-1) & MULT_71(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(51)(MULT_SIZE-1) & MULT_72(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(52)<=signed(MULT_71(52)(MULT_SIZE-1) & MULT_71(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(52)(MULT_SIZE-1) & MULT_72(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(53)<=signed(MULT_71(53)(MULT_SIZE-1) & MULT_71(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(53)(MULT_SIZE-1) & MULT_72(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(54)<=signed(MULT_71(54)(MULT_SIZE-1) & MULT_71(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(54)(MULT_SIZE-1) & MULT_72(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(55)<=signed(MULT_71(55)(MULT_SIZE-1) & MULT_71(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(55)(MULT_SIZE-1) & MULT_72(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(56)<=signed(MULT_71(56)(MULT_SIZE-1) & MULT_71(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(56)(MULT_SIZE-1) & MULT_72(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(57)<=signed(MULT_71(57)(MULT_SIZE-1) & MULT_71(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(57)(MULT_SIZE-1) & MULT_72(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(58)<=signed(MULT_71(58)(MULT_SIZE-1) & MULT_71(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(58)(MULT_SIZE-1) & MULT_72(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(59)<=signed(MULT_71(59)(MULT_SIZE-1) & MULT_71(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(59)(MULT_SIZE-1) & MULT_72(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(60)<=signed(MULT_71(60)(MULT_SIZE-1) & MULT_71(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(60)(MULT_SIZE-1) & MULT_72(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(61)<=signed(MULT_71(61)(MULT_SIZE-1) & MULT_71(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(61)(MULT_SIZE-1) & MULT_72(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(62)<=signed(MULT_71(62)(MULT_SIZE-1) & MULT_71(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(62)(MULT_SIZE-1) & MULT_72(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(63)<=signed(MULT_71(63)(MULT_SIZE-1) & MULT_71(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(63)(MULT_SIZE-1) & MULT_72(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(64)<=signed(MULT_71(64)(MULT_SIZE-1) & MULT_71(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(64)(MULT_SIZE-1) & MULT_72(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(65)<=signed(MULT_71(65)(MULT_SIZE-1) & MULT_71(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(65)(MULT_SIZE-1) & MULT_72(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(66)<=signed(MULT_71(66)(MULT_SIZE-1) & MULT_71(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(66)(MULT_SIZE-1) & MULT_72(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(67)<=signed(MULT_71(67)(MULT_SIZE-1) & MULT_71(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(67)(MULT_SIZE-1) & MULT_72(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(68)<=signed(MULT_71(68)(MULT_SIZE-1) & MULT_71(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(68)(MULT_SIZE-1) & MULT_72(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(69)<=signed(MULT_71(69)(MULT_SIZE-1) & MULT_71(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(69)(MULT_SIZE-1) & MULT_72(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(70)<=signed(MULT_71(70)(MULT_SIZE-1) & MULT_71(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(70)(MULT_SIZE-1) & MULT_72(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(71)<=signed(MULT_71(71)(MULT_SIZE-1) & MULT_71(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(71)(MULT_SIZE-1) & MULT_72(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(72)<=signed(MULT_71(72)(MULT_SIZE-1) & MULT_71(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(72)(MULT_SIZE-1) & MULT_72(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(73)<=signed(MULT_71(73)(MULT_SIZE-1) & MULT_71(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(73)(MULT_SIZE-1) & MULT_72(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(74)<=signed(MULT_71(74)(MULT_SIZE-1) & MULT_71(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(74)(MULT_SIZE-1) & MULT_72(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(75)<=signed(MULT_71(75)(MULT_SIZE-1) & MULT_71(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(75)(MULT_SIZE-1) & MULT_72(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(76)<=signed(MULT_71(76)(MULT_SIZE-1) & MULT_71(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(76)(MULT_SIZE-1) & MULT_72(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(77)<=signed(MULT_71(77)(MULT_SIZE-1) & MULT_71(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(77)(MULT_SIZE-1) & MULT_72(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(78)<=signed(MULT_71(78)(MULT_SIZE-1) & MULT_71(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(78)(MULT_SIZE-1) & MULT_72(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(79)<=signed(MULT_71(79)(MULT_SIZE-1) & MULT_71(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(79)(MULT_SIZE-1) & MULT_72(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(80)<=signed(MULT_71(80)(MULT_SIZE-1) & MULT_71(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(80)(MULT_SIZE-1) & MULT_72(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(81)<=signed(MULT_71(81)(MULT_SIZE-1) & MULT_71(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(81)(MULT_SIZE-1) & MULT_72(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(82)<=signed(MULT_71(82)(MULT_SIZE-1) & MULT_71(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(82)(MULT_SIZE-1) & MULT_72(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_36(83)<=signed(MULT_71(83)(MULT_SIZE-1) & MULT_71(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_72(83)(MULT_SIZE-1) & MULT_72(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_37(0)<=signed(MULT_73(0)(MULT_SIZE-1) & MULT_73(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(0)(MULT_SIZE-1) & MULT_74(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(1)<=signed(MULT_73(1)(MULT_SIZE-1) & MULT_73(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(1)(MULT_SIZE-1) & MULT_74(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(2)<=signed(MULT_73(2)(MULT_SIZE-1) & MULT_73(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(2)(MULT_SIZE-1) & MULT_74(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(3)<=signed(MULT_73(3)(MULT_SIZE-1) & MULT_73(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(3)(MULT_SIZE-1) & MULT_74(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(4)<=signed(MULT_73(4)(MULT_SIZE-1) & MULT_73(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(4)(MULT_SIZE-1) & MULT_74(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(5)<=signed(MULT_73(5)(MULT_SIZE-1) & MULT_73(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(5)(MULT_SIZE-1) & MULT_74(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(6)<=signed(MULT_73(6)(MULT_SIZE-1) & MULT_73(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(6)(MULT_SIZE-1) & MULT_74(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(7)<=signed(MULT_73(7)(MULT_SIZE-1) & MULT_73(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(7)(MULT_SIZE-1) & MULT_74(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(8)<=signed(MULT_73(8)(MULT_SIZE-1) & MULT_73(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(8)(MULT_SIZE-1) & MULT_74(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(9)<=signed(MULT_73(9)(MULT_SIZE-1) & MULT_73(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(9)(MULT_SIZE-1) & MULT_74(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(10)<=signed(MULT_73(10)(MULT_SIZE-1) & MULT_73(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(10)(MULT_SIZE-1) & MULT_74(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(11)<=signed(MULT_73(11)(MULT_SIZE-1) & MULT_73(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(11)(MULT_SIZE-1) & MULT_74(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(12)<=signed(MULT_73(12)(MULT_SIZE-1) & MULT_73(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(12)(MULT_SIZE-1) & MULT_74(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(13)<=signed(MULT_73(13)(MULT_SIZE-1) & MULT_73(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(13)(MULT_SIZE-1) & MULT_74(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(14)<=signed(MULT_73(14)(MULT_SIZE-1) & MULT_73(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(14)(MULT_SIZE-1) & MULT_74(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(15)<=signed(MULT_73(15)(MULT_SIZE-1) & MULT_73(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(15)(MULT_SIZE-1) & MULT_74(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(16)<=signed(MULT_73(16)(MULT_SIZE-1) & MULT_73(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(16)(MULT_SIZE-1) & MULT_74(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(17)<=signed(MULT_73(17)(MULT_SIZE-1) & MULT_73(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(17)(MULT_SIZE-1) & MULT_74(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(18)<=signed(MULT_73(18)(MULT_SIZE-1) & MULT_73(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(18)(MULT_SIZE-1) & MULT_74(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(19)<=signed(MULT_73(19)(MULT_SIZE-1) & MULT_73(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(19)(MULT_SIZE-1) & MULT_74(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(20)<=signed(MULT_73(20)(MULT_SIZE-1) & MULT_73(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(20)(MULT_SIZE-1) & MULT_74(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(21)<=signed(MULT_73(21)(MULT_SIZE-1) & MULT_73(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(21)(MULT_SIZE-1) & MULT_74(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(22)<=signed(MULT_73(22)(MULT_SIZE-1) & MULT_73(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(22)(MULT_SIZE-1) & MULT_74(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(23)<=signed(MULT_73(23)(MULT_SIZE-1) & MULT_73(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(23)(MULT_SIZE-1) & MULT_74(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(24)<=signed(MULT_73(24)(MULT_SIZE-1) & MULT_73(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(24)(MULT_SIZE-1) & MULT_74(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(25)<=signed(MULT_73(25)(MULT_SIZE-1) & MULT_73(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(25)(MULT_SIZE-1) & MULT_74(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(26)<=signed(MULT_73(26)(MULT_SIZE-1) & MULT_73(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(26)(MULT_SIZE-1) & MULT_74(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(27)<=signed(MULT_73(27)(MULT_SIZE-1) & MULT_73(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(27)(MULT_SIZE-1) & MULT_74(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(28)<=signed(MULT_73(28)(MULT_SIZE-1) & MULT_73(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(28)(MULT_SIZE-1) & MULT_74(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(29)<=signed(MULT_73(29)(MULT_SIZE-1) & MULT_73(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(29)(MULT_SIZE-1) & MULT_74(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(30)<=signed(MULT_73(30)(MULT_SIZE-1) & MULT_73(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(30)(MULT_SIZE-1) & MULT_74(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(31)<=signed(MULT_73(31)(MULT_SIZE-1) & MULT_73(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(31)(MULT_SIZE-1) & MULT_74(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(32)<=signed(MULT_73(32)(MULT_SIZE-1) & MULT_73(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(32)(MULT_SIZE-1) & MULT_74(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(33)<=signed(MULT_73(33)(MULT_SIZE-1) & MULT_73(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(33)(MULT_SIZE-1) & MULT_74(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(34)<=signed(MULT_73(34)(MULT_SIZE-1) & MULT_73(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(34)(MULT_SIZE-1) & MULT_74(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(35)<=signed(MULT_73(35)(MULT_SIZE-1) & MULT_73(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(35)(MULT_SIZE-1) & MULT_74(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(36)<=signed(MULT_73(36)(MULT_SIZE-1) & MULT_73(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(36)(MULT_SIZE-1) & MULT_74(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(37)<=signed(MULT_73(37)(MULT_SIZE-1) & MULT_73(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(37)(MULT_SIZE-1) & MULT_74(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(38)<=signed(MULT_73(38)(MULT_SIZE-1) & MULT_73(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(38)(MULT_SIZE-1) & MULT_74(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(39)<=signed(MULT_73(39)(MULT_SIZE-1) & MULT_73(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(39)(MULT_SIZE-1) & MULT_74(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(40)<=signed(MULT_73(40)(MULT_SIZE-1) & MULT_73(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(40)(MULT_SIZE-1) & MULT_74(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(41)<=signed(MULT_73(41)(MULT_SIZE-1) & MULT_73(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(41)(MULT_SIZE-1) & MULT_74(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(42)<=signed(MULT_73(42)(MULT_SIZE-1) & MULT_73(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(42)(MULT_SIZE-1) & MULT_74(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(43)<=signed(MULT_73(43)(MULT_SIZE-1) & MULT_73(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(43)(MULT_SIZE-1) & MULT_74(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(44)<=signed(MULT_73(44)(MULT_SIZE-1) & MULT_73(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(44)(MULT_SIZE-1) & MULT_74(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(45)<=signed(MULT_73(45)(MULT_SIZE-1) & MULT_73(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(45)(MULT_SIZE-1) & MULT_74(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(46)<=signed(MULT_73(46)(MULT_SIZE-1) & MULT_73(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(46)(MULT_SIZE-1) & MULT_74(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(47)<=signed(MULT_73(47)(MULT_SIZE-1) & MULT_73(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(47)(MULT_SIZE-1) & MULT_74(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(48)<=signed(MULT_73(48)(MULT_SIZE-1) & MULT_73(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(48)(MULT_SIZE-1) & MULT_74(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(49)<=signed(MULT_73(49)(MULT_SIZE-1) & MULT_73(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(49)(MULT_SIZE-1) & MULT_74(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(50)<=signed(MULT_73(50)(MULT_SIZE-1) & MULT_73(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(50)(MULT_SIZE-1) & MULT_74(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(51)<=signed(MULT_73(51)(MULT_SIZE-1) & MULT_73(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(51)(MULT_SIZE-1) & MULT_74(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(52)<=signed(MULT_73(52)(MULT_SIZE-1) & MULT_73(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(52)(MULT_SIZE-1) & MULT_74(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(53)<=signed(MULT_73(53)(MULT_SIZE-1) & MULT_73(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(53)(MULT_SIZE-1) & MULT_74(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(54)<=signed(MULT_73(54)(MULT_SIZE-1) & MULT_73(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(54)(MULT_SIZE-1) & MULT_74(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(55)<=signed(MULT_73(55)(MULT_SIZE-1) & MULT_73(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(55)(MULT_SIZE-1) & MULT_74(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(56)<=signed(MULT_73(56)(MULT_SIZE-1) & MULT_73(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(56)(MULT_SIZE-1) & MULT_74(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(57)<=signed(MULT_73(57)(MULT_SIZE-1) & MULT_73(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(57)(MULT_SIZE-1) & MULT_74(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(58)<=signed(MULT_73(58)(MULT_SIZE-1) & MULT_73(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(58)(MULT_SIZE-1) & MULT_74(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(59)<=signed(MULT_73(59)(MULT_SIZE-1) & MULT_73(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(59)(MULT_SIZE-1) & MULT_74(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(60)<=signed(MULT_73(60)(MULT_SIZE-1) & MULT_73(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(60)(MULT_SIZE-1) & MULT_74(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(61)<=signed(MULT_73(61)(MULT_SIZE-1) & MULT_73(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(61)(MULT_SIZE-1) & MULT_74(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(62)<=signed(MULT_73(62)(MULT_SIZE-1) & MULT_73(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(62)(MULT_SIZE-1) & MULT_74(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(63)<=signed(MULT_73(63)(MULT_SIZE-1) & MULT_73(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(63)(MULT_SIZE-1) & MULT_74(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(64)<=signed(MULT_73(64)(MULT_SIZE-1) & MULT_73(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(64)(MULT_SIZE-1) & MULT_74(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(65)<=signed(MULT_73(65)(MULT_SIZE-1) & MULT_73(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(65)(MULT_SIZE-1) & MULT_74(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(66)<=signed(MULT_73(66)(MULT_SIZE-1) & MULT_73(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(66)(MULT_SIZE-1) & MULT_74(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(67)<=signed(MULT_73(67)(MULT_SIZE-1) & MULT_73(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(67)(MULT_SIZE-1) & MULT_74(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(68)<=signed(MULT_73(68)(MULT_SIZE-1) & MULT_73(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(68)(MULT_SIZE-1) & MULT_74(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(69)<=signed(MULT_73(69)(MULT_SIZE-1) & MULT_73(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(69)(MULT_SIZE-1) & MULT_74(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(70)<=signed(MULT_73(70)(MULT_SIZE-1) & MULT_73(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(70)(MULT_SIZE-1) & MULT_74(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(71)<=signed(MULT_73(71)(MULT_SIZE-1) & MULT_73(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(71)(MULT_SIZE-1) & MULT_74(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(72)<=signed(MULT_73(72)(MULT_SIZE-1) & MULT_73(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(72)(MULT_SIZE-1) & MULT_74(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(73)<=signed(MULT_73(73)(MULT_SIZE-1) & MULT_73(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(73)(MULT_SIZE-1) & MULT_74(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(74)<=signed(MULT_73(74)(MULT_SIZE-1) & MULT_73(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(74)(MULT_SIZE-1) & MULT_74(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(75)<=signed(MULT_73(75)(MULT_SIZE-1) & MULT_73(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(75)(MULT_SIZE-1) & MULT_74(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(76)<=signed(MULT_73(76)(MULT_SIZE-1) & MULT_73(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(76)(MULT_SIZE-1) & MULT_74(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(77)<=signed(MULT_73(77)(MULT_SIZE-1) & MULT_73(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(77)(MULT_SIZE-1) & MULT_74(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(78)<=signed(MULT_73(78)(MULT_SIZE-1) & MULT_73(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(78)(MULT_SIZE-1) & MULT_74(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(79)<=signed(MULT_73(79)(MULT_SIZE-1) & MULT_73(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(79)(MULT_SIZE-1) & MULT_74(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(80)<=signed(MULT_73(80)(MULT_SIZE-1) & MULT_73(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(80)(MULT_SIZE-1) & MULT_74(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(81)<=signed(MULT_73(81)(MULT_SIZE-1) & MULT_73(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(81)(MULT_SIZE-1) & MULT_74(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(82)<=signed(MULT_73(82)(MULT_SIZE-1) & MULT_73(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(82)(MULT_SIZE-1) & MULT_74(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_37(83)<=signed(MULT_73(83)(MULT_SIZE-1) & MULT_73(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_74(83)(MULT_SIZE-1) & MULT_74(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_38(0)<=signed(MULT_75(0)(MULT_SIZE-1) & MULT_75(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(0)(MULT_SIZE-1) & MULT_76(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(1)<=signed(MULT_75(1)(MULT_SIZE-1) & MULT_75(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(1)(MULT_SIZE-1) & MULT_76(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(2)<=signed(MULT_75(2)(MULT_SIZE-1) & MULT_75(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(2)(MULT_SIZE-1) & MULT_76(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(3)<=signed(MULT_75(3)(MULT_SIZE-1) & MULT_75(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(3)(MULT_SIZE-1) & MULT_76(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(4)<=signed(MULT_75(4)(MULT_SIZE-1) & MULT_75(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(4)(MULT_SIZE-1) & MULT_76(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(5)<=signed(MULT_75(5)(MULT_SIZE-1) & MULT_75(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(5)(MULT_SIZE-1) & MULT_76(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(6)<=signed(MULT_75(6)(MULT_SIZE-1) & MULT_75(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(6)(MULT_SIZE-1) & MULT_76(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(7)<=signed(MULT_75(7)(MULT_SIZE-1) & MULT_75(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(7)(MULT_SIZE-1) & MULT_76(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(8)<=signed(MULT_75(8)(MULT_SIZE-1) & MULT_75(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(8)(MULT_SIZE-1) & MULT_76(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(9)<=signed(MULT_75(9)(MULT_SIZE-1) & MULT_75(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(9)(MULT_SIZE-1) & MULT_76(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(10)<=signed(MULT_75(10)(MULT_SIZE-1) & MULT_75(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(10)(MULT_SIZE-1) & MULT_76(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(11)<=signed(MULT_75(11)(MULT_SIZE-1) & MULT_75(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(11)(MULT_SIZE-1) & MULT_76(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(12)<=signed(MULT_75(12)(MULT_SIZE-1) & MULT_75(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(12)(MULT_SIZE-1) & MULT_76(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(13)<=signed(MULT_75(13)(MULT_SIZE-1) & MULT_75(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(13)(MULT_SIZE-1) & MULT_76(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(14)<=signed(MULT_75(14)(MULT_SIZE-1) & MULT_75(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(14)(MULT_SIZE-1) & MULT_76(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(15)<=signed(MULT_75(15)(MULT_SIZE-1) & MULT_75(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(15)(MULT_SIZE-1) & MULT_76(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(16)<=signed(MULT_75(16)(MULT_SIZE-1) & MULT_75(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(16)(MULT_SIZE-1) & MULT_76(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(17)<=signed(MULT_75(17)(MULT_SIZE-1) & MULT_75(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(17)(MULT_SIZE-1) & MULT_76(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(18)<=signed(MULT_75(18)(MULT_SIZE-1) & MULT_75(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(18)(MULT_SIZE-1) & MULT_76(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(19)<=signed(MULT_75(19)(MULT_SIZE-1) & MULT_75(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(19)(MULT_SIZE-1) & MULT_76(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(20)<=signed(MULT_75(20)(MULT_SIZE-1) & MULT_75(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(20)(MULT_SIZE-1) & MULT_76(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(21)<=signed(MULT_75(21)(MULT_SIZE-1) & MULT_75(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(21)(MULT_SIZE-1) & MULT_76(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(22)<=signed(MULT_75(22)(MULT_SIZE-1) & MULT_75(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(22)(MULT_SIZE-1) & MULT_76(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(23)<=signed(MULT_75(23)(MULT_SIZE-1) & MULT_75(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(23)(MULT_SIZE-1) & MULT_76(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(24)<=signed(MULT_75(24)(MULT_SIZE-1) & MULT_75(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(24)(MULT_SIZE-1) & MULT_76(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(25)<=signed(MULT_75(25)(MULT_SIZE-1) & MULT_75(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(25)(MULT_SIZE-1) & MULT_76(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(26)<=signed(MULT_75(26)(MULT_SIZE-1) & MULT_75(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(26)(MULT_SIZE-1) & MULT_76(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(27)<=signed(MULT_75(27)(MULT_SIZE-1) & MULT_75(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(27)(MULT_SIZE-1) & MULT_76(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(28)<=signed(MULT_75(28)(MULT_SIZE-1) & MULT_75(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(28)(MULT_SIZE-1) & MULT_76(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(29)<=signed(MULT_75(29)(MULT_SIZE-1) & MULT_75(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(29)(MULT_SIZE-1) & MULT_76(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(30)<=signed(MULT_75(30)(MULT_SIZE-1) & MULT_75(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(30)(MULT_SIZE-1) & MULT_76(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(31)<=signed(MULT_75(31)(MULT_SIZE-1) & MULT_75(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(31)(MULT_SIZE-1) & MULT_76(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(32)<=signed(MULT_75(32)(MULT_SIZE-1) & MULT_75(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(32)(MULT_SIZE-1) & MULT_76(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(33)<=signed(MULT_75(33)(MULT_SIZE-1) & MULT_75(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(33)(MULT_SIZE-1) & MULT_76(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(34)<=signed(MULT_75(34)(MULT_SIZE-1) & MULT_75(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(34)(MULT_SIZE-1) & MULT_76(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(35)<=signed(MULT_75(35)(MULT_SIZE-1) & MULT_75(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(35)(MULT_SIZE-1) & MULT_76(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(36)<=signed(MULT_75(36)(MULT_SIZE-1) & MULT_75(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(36)(MULT_SIZE-1) & MULT_76(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(37)<=signed(MULT_75(37)(MULT_SIZE-1) & MULT_75(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(37)(MULT_SIZE-1) & MULT_76(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(38)<=signed(MULT_75(38)(MULT_SIZE-1) & MULT_75(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(38)(MULT_SIZE-1) & MULT_76(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(39)<=signed(MULT_75(39)(MULT_SIZE-1) & MULT_75(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(39)(MULT_SIZE-1) & MULT_76(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(40)<=signed(MULT_75(40)(MULT_SIZE-1) & MULT_75(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(40)(MULT_SIZE-1) & MULT_76(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(41)<=signed(MULT_75(41)(MULT_SIZE-1) & MULT_75(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(41)(MULT_SIZE-1) & MULT_76(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(42)<=signed(MULT_75(42)(MULT_SIZE-1) & MULT_75(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(42)(MULT_SIZE-1) & MULT_76(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(43)<=signed(MULT_75(43)(MULT_SIZE-1) & MULT_75(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(43)(MULT_SIZE-1) & MULT_76(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(44)<=signed(MULT_75(44)(MULT_SIZE-1) & MULT_75(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(44)(MULT_SIZE-1) & MULT_76(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(45)<=signed(MULT_75(45)(MULT_SIZE-1) & MULT_75(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(45)(MULT_SIZE-1) & MULT_76(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(46)<=signed(MULT_75(46)(MULT_SIZE-1) & MULT_75(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(46)(MULT_SIZE-1) & MULT_76(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(47)<=signed(MULT_75(47)(MULT_SIZE-1) & MULT_75(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(47)(MULT_SIZE-1) & MULT_76(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(48)<=signed(MULT_75(48)(MULT_SIZE-1) & MULT_75(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(48)(MULT_SIZE-1) & MULT_76(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(49)<=signed(MULT_75(49)(MULT_SIZE-1) & MULT_75(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(49)(MULT_SIZE-1) & MULT_76(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(50)<=signed(MULT_75(50)(MULT_SIZE-1) & MULT_75(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(50)(MULT_SIZE-1) & MULT_76(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(51)<=signed(MULT_75(51)(MULT_SIZE-1) & MULT_75(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(51)(MULT_SIZE-1) & MULT_76(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(52)<=signed(MULT_75(52)(MULT_SIZE-1) & MULT_75(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(52)(MULT_SIZE-1) & MULT_76(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(53)<=signed(MULT_75(53)(MULT_SIZE-1) & MULT_75(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(53)(MULT_SIZE-1) & MULT_76(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(54)<=signed(MULT_75(54)(MULT_SIZE-1) & MULT_75(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(54)(MULT_SIZE-1) & MULT_76(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(55)<=signed(MULT_75(55)(MULT_SIZE-1) & MULT_75(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(55)(MULT_SIZE-1) & MULT_76(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(56)<=signed(MULT_75(56)(MULT_SIZE-1) & MULT_75(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(56)(MULT_SIZE-1) & MULT_76(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(57)<=signed(MULT_75(57)(MULT_SIZE-1) & MULT_75(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(57)(MULT_SIZE-1) & MULT_76(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(58)<=signed(MULT_75(58)(MULT_SIZE-1) & MULT_75(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(58)(MULT_SIZE-1) & MULT_76(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(59)<=signed(MULT_75(59)(MULT_SIZE-1) & MULT_75(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(59)(MULT_SIZE-1) & MULT_76(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(60)<=signed(MULT_75(60)(MULT_SIZE-1) & MULT_75(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(60)(MULT_SIZE-1) & MULT_76(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(61)<=signed(MULT_75(61)(MULT_SIZE-1) & MULT_75(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(61)(MULT_SIZE-1) & MULT_76(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(62)<=signed(MULT_75(62)(MULT_SIZE-1) & MULT_75(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(62)(MULT_SIZE-1) & MULT_76(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(63)<=signed(MULT_75(63)(MULT_SIZE-1) & MULT_75(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(63)(MULT_SIZE-1) & MULT_76(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(64)<=signed(MULT_75(64)(MULT_SIZE-1) & MULT_75(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(64)(MULT_SIZE-1) & MULT_76(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(65)<=signed(MULT_75(65)(MULT_SIZE-1) & MULT_75(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(65)(MULT_SIZE-1) & MULT_76(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(66)<=signed(MULT_75(66)(MULT_SIZE-1) & MULT_75(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(66)(MULT_SIZE-1) & MULT_76(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(67)<=signed(MULT_75(67)(MULT_SIZE-1) & MULT_75(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(67)(MULT_SIZE-1) & MULT_76(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(68)<=signed(MULT_75(68)(MULT_SIZE-1) & MULT_75(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(68)(MULT_SIZE-1) & MULT_76(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(69)<=signed(MULT_75(69)(MULT_SIZE-1) & MULT_75(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(69)(MULT_SIZE-1) & MULT_76(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(70)<=signed(MULT_75(70)(MULT_SIZE-1) & MULT_75(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(70)(MULT_SIZE-1) & MULT_76(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(71)<=signed(MULT_75(71)(MULT_SIZE-1) & MULT_75(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(71)(MULT_SIZE-1) & MULT_76(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(72)<=signed(MULT_75(72)(MULT_SIZE-1) & MULT_75(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(72)(MULT_SIZE-1) & MULT_76(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(73)<=signed(MULT_75(73)(MULT_SIZE-1) & MULT_75(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(73)(MULT_SIZE-1) & MULT_76(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(74)<=signed(MULT_75(74)(MULT_SIZE-1) & MULT_75(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(74)(MULT_SIZE-1) & MULT_76(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(75)<=signed(MULT_75(75)(MULT_SIZE-1) & MULT_75(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(75)(MULT_SIZE-1) & MULT_76(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(76)<=signed(MULT_75(76)(MULT_SIZE-1) & MULT_75(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(76)(MULT_SIZE-1) & MULT_76(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(77)<=signed(MULT_75(77)(MULT_SIZE-1) & MULT_75(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(77)(MULT_SIZE-1) & MULT_76(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(78)<=signed(MULT_75(78)(MULT_SIZE-1) & MULT_75(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(78)(MULT_SIZE-1) & MULT_76(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(79)<=signed(MULT_75(79)(MULT_SIZE-1) & MULT_75(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(79)(MULT_SIZE-1) & MULT_76(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(80)<=signed(MULT_75(80)(MULT_SIZE-1) & MULT_75(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(80)(MULT_SIZE-1) & MULT_76(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(81)<=signed(MULT_75(81)(MULT_SIZE-1) & MULT_75(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(81)(MULT_SIZE-1) & MULT_76(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(82)<=signed(MULT_75(82)(MULT_SIZE-1) & MULT_75(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(82)(MULT_SIZE-1) & MULT_76(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_38(83)<=signed(MULT_75(83)(MULT_SIZE-1) & MULT_75(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_76(83)(MULT_SIZE-1) & MULT_76(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_39(0)<=signed(MULT_77(0)(MULT_SIZE-1) & MULT_77(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(0)(MULT_SIZE-1) & MULT_78(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(1)<=signed(MULT_77(1)(MULT_SIZE-1) & MULT_77(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(1)(MULT_SIZE-1) & MULT_78(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(2)<=signed(MULT_77(2)(MULT_SIZE-1) & MULT_77(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(2)(MULT_SIZE-1) & MULT_78(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(3)<=signed(MULT_77(3)(MULT_SIZE-1) & MULT_77(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(3)(MULT_SIZE-1) & MULT_78(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(4)<=signed(MULT_77(4)(MULT_SIZE-1) & MULT_77(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(4)(MULT_SIZE-1) & MULT_78(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(5)<=signed(MULT_77(5)(MULT_SIZE-1) & MULT_77(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(5)(MULT_SIZE-1) & MULT_78(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(6)<=signed(MULT_77(6)(MULT_SIZE-1) & MULT_77(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(6)(MULT_SIZE-1) & MULT_78(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(7)<=signed(MULT_77(7)(MULT_SIZE-1) & MULT_77(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(7)(MULT_SIZE-1) & MULT_78(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(8)<=signed(MULT_77(8)(MULT_SIZE-1) & MULT_77(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(8)(MULT_SIZE-1) & MULT_78(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(9)<=signed(MULT_77(9)(MULT_SIZE-1) & MULT_77(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(9)(MULT_SIZE-1) & MULT_78(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(10)<=signed(MULT_77(10)(MULT_SIZE-1) & MULT_77(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(10)(MULT_SIZE-1) & MULT_78(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(11)<=signed(MULT_77(11)(MULT_SIZE-1) & MULT_77(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(11)(MULT_SIZE-1) & MULT_78(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(12)<=signed(MULT_77(12)(MULT_SIZE-1) & MULT_77(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(12)(MULT_SIZE-1) & MULT_78(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(13)<=signed(MULT_77(13)(MULT_SIZE-1) & MULT_77(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(13)(MULT_SIZE-1) & MULT_78(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(14)<=signed(MULT_77(14)(MULT_SIZE-1) & MULT_77(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(14)(MULT_SIZE-1) & MULT_78(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(15)<=signed(MULT_77(15)(MULT_SIZE-1) & MULT_77(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(15)(MULT_SIZE-1) & MULT_78(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(16)<=signed(MULT_77(16)(MULT_SIZE-1) & MULT_77(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(16)(MULT_SIZE-1) & MULT_78(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(17)<=signed(MULT_77(17)(MULT_SIZE-1) & MULT_77(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(17)(MULT_SIZE-1) & MULT_78(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(18)<=signed(MULT_77(18)(MULT_SIZE-1) & MULT_77(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(18)(MULT_SIZE-1) & MULT_78(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(19)<=signed(MULT_77(19)(MULT_SIZE-1) & MULT_77(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(19)(MULT_SIZE-1) & MULT_78(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(20)<=signed(MULT_77(20)(MULT_SIZE-1) & MULT_77(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(20)(MULT_SIZE-1) & MULT_78(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(21)<=signed(MULT_77(21)(MULT_SIZE-1) & MULT_77(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(21)(MULT_SIZE-1) & MULT_78(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(22)<=signed(MULT_77(22)(MULT_SIZE-1) & MULT_77(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(22)(MULT_SIZE-1) & MULT_78(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(23)<=signed(MULT_77(23)(MULT_SIZE-1) & MULT_77(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(23)(MULT_SIZE-1) & MULT_78(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(24)<=signed(MULT_77(24)(MULT_SIZE-1) & MULT_77(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(24)(MULT_SIZE-1) & MULT_78(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(25)<=signed(MULT_77(25)(MULT_SIZE-1) & MULT_77(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(25)(MULT_SIZE-1) & MULT_78(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(26)<=signed(MULT_77(26)(MULT_SIZE-1) & MULT_77(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(26)(MULT_SIZE-1) & MULT_78(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(27)<=signed(MULT_77(27)(MULT_SIZE-1) & MULT_77(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(27)(MULT_SIZE-1) & MULT_78(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(28)<=signed(MULT_77(28)(MULT_SIZE-1) & MULT_77(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(28)(MULT_SIZE-1) & MULT_78(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(29)<=signed(MULT_77(29)(MULT_SIZE-1) & MULT_77(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(29)(MULT_SIZE-1) & MULT_78(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(30)<=signed(MULT_77(30)(MULT_SIZE-1) & MULT_77(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(30)(MULT_SIZE-1) & MULT_78(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(31)<=signed(MULT_77(31)(MULT_SIZE-1) & MULT_77(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(31)(MULT_SIZE-1) & MULT_78(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(32)<=signed(MULT_77(32)(MULT_SIZE-1) & MULT_77(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(32)(MULT_SIZE-1) & MULT_78(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(33)<=signed(MULT_77(33)(MULT_SIZE-1) & MULT_77(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(33)(MULT_SIZE-1) & MULT_78(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(34)<=signed(MULT_77(34)(MULT_SIZE-1) & MULT_77(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(34)(MULT_SIZE-1) & MULT_78(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(35)<=signed(MULT_77(35)(MULT_SIZE-1) & MULT_77(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(35)(MULT_SIZE-1) & MULT_78(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(36)<=signed(MULT_77(36)(MULT_SIZE-1) & MULT_77(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(36)(MULT_SIZE-1) & MULT_78(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(37)<=signed(MULT_77(37)(MULT_SIZE-1) & MULT_77(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(37)(MULT_SIZE-1) & MULT_78(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(38)<=signed(MULT_77(38)(MULT_SIZE-1) & MULT_77(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(38)(MULT_SIZE-1) & MULT_78(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(39)<=signed(MULT_77(39)(MULT_SIZE-1) & MULT_77(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(39)(MULT_SIZE-1) & MULT_78(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(40)<=signed(MULT_77(40)(MULT_SIZE-1) & MULT_77(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(40)(MULT_SIZE-1) & MULT_78(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(41)<=signed(MULT_77(41)(MULT_SIZE-1) & MULT_77(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(41)(MULT_SIZE-1) & MULT_78(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(42)<=signed(MULT_77(42)(MULT_SIZE-1) & MULT_77(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(42)(MULT_SIZE-1) & MULT_78(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(43)<=signed(MULT_77(43)(MULT_SIZE-1) & MULT_77(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(43)(MULT_SIZE-1) & MULT_78(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(44)<=signed(MULT_77(44)(MULT_SIZE-1) & MULT_77(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(44)(MULT_SIZE-1) & MULT_78(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(45)<=signed(MULT_77(45)(MULT_SIZE-1) & MULT_77(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(45)(MULT_SIZE-1) & MULT_78(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(46)<=signed(MULT_77(46)(MULT_SIZE-1) & MULT_77(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(46)(MULT_SIZE-1) & MULT_78(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(47)<=signed(MULT_77(47)(MULT_SIZE-1) & MULT_77(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(47)(MULT_SIZE-1) & MULT_78(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(48)<=signed(MULT_77(48)(MULT_SIZE-1) & MULT_77(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(48)(MULT_SIZE-1) & MULT_78(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(49)<=signed(MULT_77(49)(MULT_SIZE-1) & MULT_77(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(49)(MULT_SIZE-1) & MULT_78(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(50)<=signed(MULT_77(50)(MULT_SIZE-1) & MULT_77(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(50)(MULT_SIZE-1) & MULT_78(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(51)<=signed(MULT_77(51)(MULT_SIZE-1) & MULT_77(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(51)(MULT_SIZE-1) & MULT_78(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(52)<=signed(MULT_77(52)(MULT_SIZE-1) & MULT_77(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(52)(MULT_SIZE-1) & MULT_78(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(53)<=signed(MULT_77(53)(MULT_SIZE-1) & MULT_77(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(53)(MULT_SIZE-1) & MULT_78(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(54)<=signed(MULT_77(54)(MULT_SIZE-1) & MULT_77(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(54)(MULT_SIZE-1) & MULT_78(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(55)<=signed(MULT_77(55)(MULT_SIZE-1) & MULT_77(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(55)(MULT_SIZE-1) & MULT_78(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(56)<=signed(MULT_77(56)(MULT_SIZE-1) & MULT_77(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(56)(MULT_SIZE-1) & MULT_78(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(57)<=signed(MULT_77(57)(MULT_SIZE-1) & MULT_77(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(57)(MULT_SIZE-1) & MULT_78(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(58)<=signed(MULT_77(58)(MULT_SIZE-1) & MULT_77(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(58)(MULT_SIZE-1) & MULT_78(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(59)<=signed(MULT_77(59)(MULT_SIZE-1) & MULT_77(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(59)(MULT_SIZE-1) & MULT_78(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(60)<=signed(MULT_77(60)(MULT_SIZE-1) & MULT_77(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(60)(MULT_SIZE-1) & MULT_78(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(61)<=signed(MULT_77(61)(MULT_SIZE-1) & MULT_77(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(61)(MULT_SIZE-1) & MULT_78(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(62)<=signed(MULT_77(62)(MULT_SIZE-1) & MULT_77(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(62)(MULT_SIZE-1) & MULT_78(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(63)<=signed(MULT_77(63)(MULT_SIZE-1) & MULT_77(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(63)(MULT_SIZE-1) & MULT_78(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(64)<=signed(MULT_77(64)(MULT_SIZE-1) & MULT_77(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(64)(MULT_SIZE-1) & MULT_78(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(65)<=signed(MULT_77(65)(MULT_SIZE-1) & MULT_77(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(65)(MULT_SIZE-1) & MULT_78(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(66)<=signed(MULT_77(66)(MULT_SIZE-1) & MULT_77(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(66)(MULT_SIZE-1) & MULT_78(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(67)<=signed(MULT_77(67)(MULT_SIZE-1) & MULT_77(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(67)(MULT_SIZE-1) & MULT_78(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(68)<=signed(MULT_77(68)(MULT_SIZE-1) & MULT_77(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(68)(MULT_SIZE-1) & MULT_78(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(69)<=signed(MULT_77(69)(MULT_SIZE-1) & MULT_77(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(69)(MULT_SIZE-1) & MULT_78(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(70)<=signed(MULT_77(70)(MULT_SIZE-1) & MULT_77(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(70)(MULT_SIZE-1) & MULT_78(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(71)<=signed(MULT_77(71)(MULT_SIZE-1) & MULT_77(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(71)(MULT_SIZE-1) & MULT_78(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(72)<=signed(MULT_77(72)(MULT_SIZE-1) & MULT_77(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(72)(MULT_SIZE-1) & MULT_78(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(73)<=signed(MULT_77(73)(MULT_SIZE-1) & MULT_77(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(73)(MULT_SIZE-1) & MULT_78(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(74)<=signed(MULT_77(74)(MULT_SIZE-1) & MULT_77(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(74)(MULT_SIZE-1) & MULT_78(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(75)<=signed(MULT_77(75)(MULT_SIZE-1) & MULT_77(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(75)(MULT_SIZE-1) & MULT_78(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(76)<=signed(MULT_77(76)(MULT_SIZE-1) & MULT_77(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(76)(MULT_SIZE-1) & MULT_78(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(77)<=signed(MULT_77(77)(MULT_SIZE-1) & MULT_77(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(77)(MULT_SIZE-1) & MULT_78(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(78)<=signed(MULT_77(78)(MULT_SIZE-1) & MULT_77(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(78)(MULT_SIZE-1) & MULT_78(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(79)<=signed(MULT_77(79)(MULT_SIZE-1) & MULT_77(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(79)(MULT_SIZE-1) & MULT_78(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(80)<=signed(MULT_77(80)(MULT_SIZE-1) & MULT_77(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(80)(MULT_SIZE-1) & MULT_78(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(81)<=signed(MULT_77(81)(MULT_SIZE-1) & MULT_77(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(81)(MULT_SIZE-1) & MULT_78(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(82)<=signed(MULT_77(82)(MULT_SIZE-1) & MULT_77(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(82)(MULT_SIZE-1) & MULT_78(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_39(83)<=signed(MULT_77(83)(MULT_SIZE-1) & MULT_77(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_78(83)(MULT_SIZE-1) & MULT_78(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_40(0)<=signed(MULT_79(0)(MULT_SIZE-1) & MULT_79(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(0)(MULT_SIZE-1) & MULT_80(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(1)<=signed(MULT_79(1)(MULT_SIZE-1) & MULT_79(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(1)(MULT_SIZE-1) & MULT_80(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(2)<=signed(MULT_79(2)(MULT_SIZE-1) & MULT_79(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(2)(MULT_SIZE-1) & MULT_80(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(3)<=signed(MULT_79(3)(MULT_SIZE-1) & MULT_79(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(3)(MULT_SIZE-1) & MULT_80(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(4)<=signed(MULT_79(4)(MULT_SIZE-1) & MULT_79(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(4)(MULT_SIZE-1) & MULT_80(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(5)<=signed(MULT_79(5)(MULT_SIZE-1) & MULT_79(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(5)(MULT_SIZE-1) & MULT_80(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(6)<=signed(MULT_79(6)(MULT_SIZE-1) & MULT_79(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(6)(MULT_SIZE-1) & MULT_80(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(7)<=signed(MULT_79(7)(MULT_SIZE-1) & MULT_79(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(7)(MULT_SIZE-1) & MULT_80(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(8)<=signed(MULT_79(8)(MULT_SIZE-1) & MULT_79(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(8)(MULT_SIZE-1) & MULT_80(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(9)<=signed(MULT_79(9)(MULT_SIZE-1) & MULT_79(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(9)(MULT_SIZE-1) & MULT_80(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(10)<=signed(MULT_79(10)(MULT_SIZE-1) & MULT_79(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(10)(MULT_SIZE-1) & MULT_80(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(11)<=signed(MULT_79(11)(MULT_SIZE-1) & MULT_79(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(11)(MULT_SIZE-1) & MULT_80(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(12)<=signed(MULT_79(12)(MULT_SIZE-1) & MULT_79(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(12)(MULT_SIZE-1) & MULT_80(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(13)<=signed(MULT_79(13)(MULT_SIZE-1) & MULT_79(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(13)(MULT_SIZE-1) & MULT_80(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(14)<=signed(MULT_79(14)(MULT_SIZE-1) & MULT_79(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(14)(MULT_SIZE-1) & MULT_80(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(15)<=signed(MULT_79(15)(MULT_SIZE-1) & MULT_79(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(15)(MULT_SIZE-1) & MULT_80(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(16)<=signed(MULT_79(16)(MULT_SIZE-1) & MULT_79(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(16)(MULT_SIZE-1) & MULT_80(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(17)<=signed(MULT_79(17)(MULT_SIZE-1) & MULT_79(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(17)(MULT_SIZE-1) & MULT_80(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(18)<=signed(MULT_79(18)(MULT_SIZE-1) & MULT_79(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(18)(MULT_SIZE-1) & MULT_80(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(19)<=signed(MULT_79(19)(MULT_SIZE-1) & MULT_79(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(19)(MULT_SIZE-1) & MULT_80(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(20)<=signed(MULT_79(20)(MULT_SIZE-1) & MULT_79(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(20)(MULT_SIZE-1) & MULT_80(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(21)<=signed(MULT_79(21)(MULT_SIZE-1) & MULT_79(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(21)(MULT_SIZE-1) & MULT_80(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(22)<=signed(MULT_79(22)(MULT_SIZE-1) & MULT_79(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(22)(MULT_SIZE-1) & MULT_80(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(23)<=signed(MULT_79(23)(MULT_SIZE-1) & MULT_79(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(23)(MULT_SIZE-1) & MULT_80(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(24)<=signed(MULT_79(24)(MULT_SIZE-1) & MULT_79(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(24)(MULT_SIZE-1) & MULT_80(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(25)<=signed(MULT_79(25)(MULT_SIZE-1) & MULT_79(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(25)(MULT_SIZE-1) & MULT_80(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(26)<=signed(MULT_79(26)(MULT_SIZE-1) & MULT_79(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(26)(MULT_SIZE-1) & MULT_80(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(27)<=signed(MULT_79(27)(MULT_SIZE-1) & MULT_79(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(27)(MULT_SIZE-1) & MULT_80(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(28)<=signed(MULT_79(28)(MULT_SIZE-1) & MULT_79(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(28)(MULT_SIZE-1) & MULT_80(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(29)<=signed(MULT_79(29)(MULT_SIZE-1) & MULT_79(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(29)(MULT_SIZE-1) & MULT_80(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(30)<=signed(MULT_79(30)(MULT_SIZE-1) & MULT_79(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(30)(MULT_SIZE-1) & MULT_80(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(31)<=signed(MULT_79(31)(MULT_SIZE-1) & MULT_79(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(31)(MULT_SIZE-1) & MULT_80(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(32)<=signed(MULT_79(32)(MULT_SIZE-1) & MULT_79(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(32)(MULT_SIZE-1) & MULT_80(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(33)<=signed(MULT_79(33)(MULT_SIZE-1) & MULT_79(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(33)(MULT_SIZE-1) & MULT_80(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(34)<=signed(MULT_79(34)(MULT_SIZE-1) & MULT_79(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(34)(MULT_SIZE-1) & MULT_80(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(35)<=signed(MULT_79(35)(MULT_SIZE-1) & MULT_79(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(35)(MULT_SIZE-1) & MULT_80(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(36)<=signed(MULT_79(36)(MULT_SIZE-1) & MULT_79(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(36)(MULT_SIZE-1) & MULT_80(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(37)<=signed(MULT_79(37)(MULT_SIZE-1) & MULT_79(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(37)(MULT_SIZE-1) & MULT_80(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(38)<=signed(MULT_79(38)(MULT_SIZE-1) & MULT_79(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(38)(MULT_SIZE-1) & MULT_80(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(39)<=signed(MULT_79(39)(MULT_SIZE-1) & MULT_79(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(39)(MULT_SIZE-1) & MULT_80(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(40)<=signed(MULT_79(40)(MULT_SIZE-1) & MULT_79(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(40)(MULT_SIZE-1) & MULT_80(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(41)<=signed(MULT_79(41)(MULT_SIZE-1) & MULT_79(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(41)(MULT_SIZE-1) & MULT_80(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(42)<=signed(MULT_79(42)(MULT_SIZE-1) & MULT_79(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(42)(MULT_SIZE-1) & MULT_80(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(43)<=signed(MULT_79(43)(MULT_SIZE-1) & MULT_79(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(43)(MULT_SIZE-1) & MULT_80(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(44)<=signed(MULT_79(44)(MULT_SIZE-1) & MULT_79(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(44)(MULT_SIZE-1) & MULT_80(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(45)<=signed(MULT_79(45)(MULT_SIZE-1) & MULT_79(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(45)(MULT_SIZE-1) & MULT_80(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(46)<=signed(MULT_79(46)(MULT_SIZE-1) & MULT_79(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(46)(MULT_SIZE-1) & MULT_80(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(47)<=signed(MULT_79(47)(MULT_SIZE-1) & MULT_79(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(47)(MULT_SIZE-1) & MULT_80(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(48)<=signed(MULT_79(48)(MULT_SIZE-1) & MULT_79(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(48)(MULT_SIZE-1) & MULT_80(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(49)<=signed(MULT_79(49)(MULT_SIZE-1) & MULT_79(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(49)(MULT_SIZE-1) & MULT_80(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(50)<=signed(MULT_79(50)(MULT_SIZE-1) & MULT_79(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(50)(MULT_SIZE-1) & MULT_80(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(51)<=signed(MULT_79(51)(MULT_SIZE-1) & MULT_79(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(51)(MULT_SIZE-1) & MULT_80(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(52)<=signed(MULT_79(52)(MULT_SIZE-1) & MULT_79(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(52)(MULT_SIZE-1) & MULT_80(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(53)<=signed(MULT_79(53)(MULT_SIZE-1) & MULT_79(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(53)(MULT_SIZE-1) & MULT_80(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(54)<=signed(MULT_79(54)(MULT_SIZE-1) & MULT_79(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(54)(MULT_SIZE-1) & MULT_80(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(55)<=signed(MULT_79(55)(MULT_SIZE-1) & MULT_79(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(55)(MULT_SIZE-1) & MULT_80(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(56)<=signed(MULT_79(56)(MULT_SIZE-1) & MULT_79(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(56)(MULT_SIZE-1) & MULT_80(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(57)<=signed(MULT_79(57)(MULT_SIZE-1) & MULT_79(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(57)(MULT_SIZE-1) & MULT_80(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(58)<=signed(MULT_79(58)(MULT_SIZE-1) & MULT_79(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(58)(MULT_SIZE-1) & MULT_80(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(59)<=signed(MULT_79(59)(MULT_SIZE-1) & MULT_79(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(59)(MULT_SIZE-1) & MULT_80(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(60)<=signed(MULT_79(60)(MULT_SIZE-1) & MULT_79(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(60)(MULT_SIZE-1) & MULT_80(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(61)<=signed(MULT_79(61)(MULT_SIZE-1) & MULT_79(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(61)(MULT_SIZE-1) & MULT_80(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(62)<=signed(MULT_79(62)(MULT_SIZE-1) & MULT_79(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(62)(MULT_SIZE-1) & MULT_80(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(63)<=signed(MULT_79(63)(MULT_SIZE-1) & MULT_79(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(63)(MULT_SIZE-1) & MULT_80(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(64)<=signed(MULT_79(64)(MULT_SIZE-1) & MULT_79(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(64)(MULT_SIZE-1) & MULT_80(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(65)<=signed(MULT_79(65)(MULT_SIZE-1) & MULT_79(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(65)(MULT_SIZE-1) & MULT_80(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(66)<=signed(MULT_79(66)(MULT_SIZE-1) & MULT_79(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(66)(MULT_SIZE-1) & MULT_80(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(67)<=signed(MULT_79(67)(MULT_SIZE-1) & MULT_79(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(67)(MULT_SIZE-1) & MULT_80(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(68)<=signed(MULT_79(68)(MULT_SIZE-1) & MULT_79(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(68)(MULT_SIZE-1) & MULT_80(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(69)<=signed(MULT_79(69)(MULT_SIZE-1) & MULT_79(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(69)(MULT_SIZE-1) & MULT_80(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(70)<=signed(MULT_79(70)(MULT_SIZE-1) & MULT_79(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(70)(MULT_SIZE-1) & MULT_80(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(71)<=signed(MULT_79(71)(MULT_SIZE-1) & MULT_79(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(71)(MULT_SIZE-1) & MULT_80(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(72)<=signed(MULT_79(72)(MULT_SIZE-1) & MULT_79(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(72)(MULT_SIZE-1) & MULT_80(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(73)<=signed(MULT_79(73)(MULT_SIZE-1) & MULT_79(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(73)(MULT_SIZE-1) & MULT_80(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(74)<=signed(MULT_79(74)(MULT_SIZE-1) & MULT_79(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(74)(MULT_SIZE-1) & MULT_80(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(75)<=signed(MULT_79(75)(MULT_SIZE-1) & MULT_79(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(75)(MULT_SIZE-1) & MULT_80(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(76)<=signed(MULT_79(76)(MULT_SIZE-1) & MULT_79(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(76)(MULT_SIZE-1) & MULT_80(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(77)<=signed(MULT_79(77)(MULT_SIZE-1) & MULT_79(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(77)(MULT_SIZE-1) & MULT_80(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(78)<=signed(MULT_79(78)(MULT_SIZE-1) & MULT_79(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(78)(MULT_SIZE-1) & MULT_80(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(79)<=signed(MULT_79(79)(MULT_SIZE-1) & MULT_79(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(79)(MULT_SIZE-1) & MULT_80(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(80)<=signed(MULT_79(80)(MULT_SIZE-1) & MULT_79(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(80)(MULT_SIZE-1) & MULT_80(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(81)<=signed(MULT_79(81)(MULT_SIZE-1) & MULT_79(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(81)(MULT_SIZE-1) & MULT_80(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(82)<=signed(MULT_79(82)(MULT_SIZE-1) & MULT_79(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(82)(MULT_SIZE-1) & MULT_80(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_40(83)<=signed(MULT_79(83)(MULT_SIZE-1) & MULT_79(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_80(83)(MULT_SIZE-1) & MULT_80(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_41(0)<=signed(MULT_81(0)(MULT_SIZE-1) & MULT_81(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(0)(MULT_SIZE-1) & MULT_82(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(1)<=signed(MULT_81(1)(MULT_SIZE-1) & MULT_81(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(1)(MULT_SIZE-1) & MULT_82(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(2)<=signed(MULT_81(2)(MULT_SIZE-1) & MULT_81(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(2)(MULT_SIZE-1) & MULT_82(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(3)<=signed(MULT_81(3)(MULT_SIZE-1) & MULT_81(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(3)(MULT_SIZE-1) & MULT_82(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(4)<=signed(MULT_81(4)(MULT_SIZE-1) & MULT_81(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(4)(MULT_SIZE-1) & MULT_82(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(5)<=signed(MULT_81(5)(MULT_SIZE-1) & MULT_81(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(5)(MULT_SIZE-1) & MULT_82(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(6)<=signed(MULT_81(6)(MULT_SIZE-1) & MULT_81(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(6)(MULT_SIZE-1) & MULT_82(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(7)<=signed(MULT_81(7)(MULT_SIZE-1) & MULT_81(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(7)(MULT_SIZE-1) & MULT_82(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(8)<=signed(MULT_81(8)(MULT_SIZE-1) & MULT_81(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(8)(MULT_SIZE-1) & MULT_82(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(9)<=signed(MULT_81(9)(MULT_SIZE-1) & MULT_81(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(9)(MULT_SIZE-1) & MULT_82(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(10)<=signed(MULT_81(10)(MULT_SIZE-1) & MULT_81(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(10)(MULT_SIZE-1) & MULT_82(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(11)<=signed(MULT_81(11)(MULT_SIZE-1) & MULT_81(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(11)(MULT_SIZE-1) & MULT_82(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(12)<=signed(MULT_81(12)(MULT_SIZE-1) & MULT_81(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(12)(MULT_SIZE-1) & MULT_82(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(13)<=signed(MULT_81(13)(MULT_SIZE-1) & MULT_81(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(13)(MULT_SIZE-1) & MULT_82(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(14)<=signed(MULT_81(14)(MULT_SIZE-1) & MULT_81(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(14)(MULT_SIZE-1) & MULT_82(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(15)<=signed(MULT_81(15)(MULT_SIZE-1) & MULT_81(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(15)(MULT_SIZE-1) & MULT_82(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(16)<=signed(MULT_81(16)(MULT_SIZE-1) & MULT_81(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(16)(MULT_SIZE-1) & MULT_82(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(17)<=signed(MULT_81(17)(MULT_SIZE-1) & MULT_81(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(17)(MULT_SIZE-1) & MULT_82(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(18)<=signed(MULT_81(18)(MULT_SIZE-1) & MULT_81(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(18)(MULT_SIZE-1) & MULT_82(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(19)<=signed(MULT_81(19)(MULT_SIZE-1) & MULT_81(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(19)(MULT_SIZE-1) & MULT_82(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(20)<=signed(MULT_81(20)(MULT_SIZE-1) & MULT_81(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(20)(MULT_SIZE-1) & MULT_82(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(21)<=signed(MULT_81(21)(MULT_SIZE-1) & MULT_81(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(21)(MULT_SIZE-1) & MULT_82(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(22)<=signed(MULT_81(22)(MULT_SIZE-1) & MULT_81(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(22)(MULT_SIZE-1) & MULT_82(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(23)<=signed(MULT_81(23)(MULT_SIZE-1) & MULT_81(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(23)(MULT_SIZE-1) & MULT_82(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(24)<=signed(MULT_81(24)(MULT_SIZE-1) & MULT_81(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(24)(MULT_SIZE-1) & MULT_82(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(25)<=signed(MULT_81(25)(MULT_SIZE-1) & MULT_81(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(25)(MULT_SIZE-1) & MULT_82(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(26)<=signed(MULT_81(26)(MULT_SIZE-1) & MULT_81(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(26)(MULT_SIZE-1) & MULT_82(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(27)<=signed(MULT_81(27)(MULT_SIZE-1) & MULT_81(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(27)(MULT_SIZE-1) & MULT_82(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(28)<=signed(MULT_81(28)(MULT_SIZE-1) & MULT_81(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(28)(MULT_SIZE-1) & MULT_82(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(29)<=signed(MULT_81(29)(MULT_SIZE-1) & MULT_81(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(29)(MULT_SIZE-1) & MULT_82(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(30)<=signed(MULT_81(30)(MULT_SIZE-1) & MULT_81(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(30)(MULT_SIZE-1) & MULT_82(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(31)<=signed(MULT_81(31)(MULT_SIZE-1) & MULT_81(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(31)(MULT_SIZE-1) & MULT_82(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(32)<=signed(MULT_81(32)(MULT_SIZE-1) & MULT_81(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(32)(MULT_SIZE-1) & MULT_82(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(33)<=signed(MULT_81(33)(MULT_SIZE-1) & MULT_81(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(33)(MULT_SIZE-1) & MULT_82(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(34)<=signed(MULT_81(34)(MULT_SIZE-1) & MULT_81(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(34)(MULT_SIZE-1) & MULT_82(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(35)<=signed(MULT_81(35)(MULT_SIZE-1) & MULT_81(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(35)(MULT_SIZE-1) & MULT_82(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(36)<=signed(MULT_81(36)(MULT_SIZE-1) & MULT_81(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(36)(MULT_SIZE-1) & MULT_82(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(37)<=signed(MULT_81(37)(MULT_SIZE-1) & MULT_81(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(37)(MULT_SIZE-1) & MULT_82(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(38)<=signed(MULT_81(38)(MULT_SIZE-1) & MULT_81(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(38)(MULT_SIZE-1) & MULT_82(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(39)<=signed(MULT_81(39)(MULT_SIZE-1) & MULT_81(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(39)(MULT_SIZE-1) & MULT_82(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(40)<=signed(MULT_81(40)(MULT_SIZE-1) & MULT_81(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(40)(MULT_SIZE-1) & MULT_82(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(41)<=signed(MULT_81(41)(MULT_SIZE-1) & MULT_81(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(41)(MULT_SIZE-1) & MULT_82(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(42)<=signed(MULT_81(42)(MULT_SIZE-1) & MULT_81(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(42)(MULT_SIZE-1) & MULT_82(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(43)<=signed(MULT_81(43)(MULT_SIZE-1) & MULT_81(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(43)(MULT_SIZE-1) & MULT_82(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(44)<=signed(MULT_81(44)(MULT_SIZE-1) & MULT_81(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(44)(MULT_SIZE-1) & MULT_82(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(45)<=signed(MULT_81(45)(MULT_SIZE-1) & MULT_81(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(45)(MULT_SIZE-1) & MULT_82(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(46)<=signed(MULT_81(46)(MULT_SIZE-1) & MULT_81(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(46)(MULT_SIZE-1) & MULT_82(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(47)<=signed(MULT_81(47)(MULT_SIZE-1) & MULT_81(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(47)(MULT_SIZE-1) & MULT_82(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(48)<=signed(MULT_81(48)(MULT_SIZE-1) & MULT_81(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(48)(MULT_SIZE-1) & MULT_82(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(49)<=signed(MULT_81(49)(MULT_SIZE-1) & MULT_81(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(49)(MULT_SIZE-1) & MULT_82(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(50)<=signed(MULT_81(50)(MULT_SIZE-1) & MULT_81(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(50)(MULT_SIZE-1) & MULT_82(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(51)<=signed(MULT_81(51)(MULT_SIZE-1) & MULT_81(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(51)(MULT_SIZE-1) & MULT_82(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(52)<=signed(MULT_81(52)(MULT_SIZE-1) & MULT_81(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(52)(MULT_SIZE-1) & MULT_82(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(53)<=signed(MULT_81(53)(MULT_SIZE-1) & MULT_81(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(53)(MULT_SIZE-1) & MULT_82(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(54)<=signed(MULT_81(54)(MULT_SIZE-1) & MULT_81(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(54)(MULT_SIZE-1) & MULT_82(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(55)<=signed(MULT_81(55)(MULT_SIZE-1) & MULT_81(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(55)(MULT_SIZE-1) & MULT_82(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(56)<=signed(MULT_81(56)(MULT_SIZE-1) & MULT_81(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(56)(MULT_SIZE-1) & MULT_82(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(57)<=signed(MULT_81(57)(MULT_SIZE-1) & MULT_81(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(57)(MULT_SIZE-1) & MULT_82(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(58)<=signed(MULT_81(58)(MULT_SIZE-1) & MULT_81(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(58)(MULT_SIZE-1) & MULT_82(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(59)<=signed(MULT_81(59)(MULT_SIZE-1) & MULT_81(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(59)(MULT_SIZE-1) & MULT_82(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(60)<=signed(MULT_81(60)(MULT_SIZE-1) & MULT_81(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(60)(MULT_SIZE-1) & MULT_82(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(61)<=signed(MULT_81(61)(MULT_SIZE-1) & MULT_81(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(61)(MULT_SIZE-1) & MULT_82(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(62)<=signed(MULT_81(62)(MULT_SIZE-1) & MULT_81(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(62)(MULT_SIZE-1) & MULT_82(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(63)<=signed(MULT_81(63)(MULT_SIZE-1) & MULT_81(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(63)(MULT_SIZE-1) & MULT_82(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(64)<=signed(MULT_81(64)(MULT_SIZE-1) & MULT_81(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(64)(MULT_SIZE-1) & MULT_82(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(65)<=signed(MULT_81(65)(MULT_SIZE-1) & MULT_81(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(65)(MULT_SIZE-1) & MULT_82(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(66)<=signed(MULT_81(66)(MULT_SIZE-1) & MULT_81(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(66)(MULT_SIZE-1) & MULT_82(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(67)<=signed(MULT_81(67)(MULT_SIZE-1) & MULT_81(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(67)(MULT_SIZE-1) & MULT_82(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(68)<=signed(MULT_81(68)(MULT_SIZE-1) & MULT_81(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(68)(MULT_SIZE-1) & MULT_82(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(69)<=signed(MULT_81(69)(MULT_SIZE-1) & MULT_81(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(69)(MULT_SIZE-1) & MULT_82(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(70)<=signed(MULT_81(70)(MULT_SIZE-1) & MULT_81(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(70)(MULT_SIZE-1) & MULT_82(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(71)<=signed(MULT_81(71)(MULT_SIZE-1) & MULT_81(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(71)(MULT_SIZE-1) & MULT_82(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(72)<=signed(MULT_81(72)(MULT_SIZE-1) & MULT_81(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(72)(MULT_SIZE-1) & MULT_82(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(73)<=signed(MULT_81(73)(MULT_SIZE-1) & MULT_81(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(73)(MULT_SIZE-1) & MULT_82(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(74)<=signed(MULT_81(74)(MULT_SIZE-1) & MULT_81(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(74)(MULT_SIZE-1) & MULT_82(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(75)<=signed(MULT_81(75)(MULT_SIZE-1) & MULT_81(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(75)(MULT_SIZE-1) & MULT_82(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(76)<=signed(MULT_81(76)(MULT_SIZE-1) & MULT_81(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(76)(MULT_SIZE-1) & MULT_82(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(77)<=signed(MULT_81(77)(MULT_SIZE-1) & MULT_81(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(77)(MULT_SIZE-1) & MULT_82(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(78)<=signed(MULT_81(78)(MULT_SIZE-1) & MULT_81(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(78)(MULT_SIZE-1) & MULT_82(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(79)<=signed(MULT_81(79)(MULT_SIZE-1) & MULT_81(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(79)(MULT_SIZE-1) & MULT_82(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(80)<=signed(MULT_81(80)(MULT_SIZE-1) & MULT_81(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(80)(MULT_SIZE-1) & MULT_82(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(81)<=signed(MULT_81(81)(MULT_SIZE-1) & MULT_81(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(81)(MULT_SIZE-1) & MULT_82(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(82)<=signed(MULT_81(82)(MULT_SIZE-1) & MULT_81(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(82)(MULT_SIZE-1) & MULT_82(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_41(83)<=signed(MULT_81(83)(MULT_SIZE-1) & MULT_81(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_82(83)(MULT_SIZE-1) & MULT_82(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_42(0)<=signed(MULT_83(0)(MULT_SIZE-1) & MULT_83(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(0)(MULT_SIZE-1) & MULT_84(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(1)<=signed(MULT_83(1)(MULT_SIZE-1) & MULT_83(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(1)(MULT_SIZE-1) & MULT_84(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(2)<=signed(MULT_83(2)(MULT_SIZE-1) & MULT_83(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(2)(MULT_SIZE-1) & MULT_84(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(3)<=signed(MULT_83(3)(MULT_SIZE-1) & MULT_83(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(3)(MULT_SIZE-1) & MULT_84(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(4)<=signed(MULT_83(4)(MULT_SIZE-1) & MULT_83(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(4)(MULT_SIZE-1) & MULT_84(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(5)<=signed(MULT_83(5)(MULT_SIZE-1) & MULT_83(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(5)(MULT_SIZE-1) & MULT_84(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(6)<=signed(MULT_83(6)(MULT_SIZE-1) & MULT_83(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(6)(MULT_SIZE-1) & MULT_84(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(7)<=signed(MULT_83(7)(MULT_SIZE-1) & MULT_83(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(7)(MULT_SIZE-1) & MULT_84(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(8)<=signed(MULT_83(8)(MULT_SIZE-1) & MULT_83(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(8)(MULT_SIZE-1) & MULT_84(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(9)<=signed(MULT_83(9)(MULT_SIZE-1) & MULT_83(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(9)(MULT_SIZE-1) & MULT_84(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(10)<=signed(MULT_83(10)(MULT_SIZE-1) & MULT_83(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(10)(MULT_SIZE-1) & MULT_84(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(11)<=signed(MULT_83(11)(MULT_SIZE-1) & MULT_83(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(11)(MULT_SIZE-1) & MULT_84(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(12)<=signed(MULT_83(12)(MULT_SIZE-1) & MULT_83(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(12)(MULT_SIZE-1) & MULT_84(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(13)<=signed(MULT_83(13)(MULT_SIZE-1) & MULT_83(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(13)(MULT_SIZE-1) & MULT_84(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(14)<=signed(MULT_83(14)(MULT_SIZE-1) & MULT_83(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(14)(MULT_SIZE-1) & MULT_84(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(15)<=signed(MULT_83(15)(MULT_SIZE-1) & MULT_83(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(15)(MULT_SIZE-1) & MULT_84(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(16)<=signed(MULT_83(16)(MULT_SIZE-1) & MULT_83(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(16)(MULT_SIZE-1) & MULT_84(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(17)<=signed(MULT_83(17)(MULT_SIZE-1) & MULT_83(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(17)(MULT_SIZE-1) & MULT_84(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(18)<=signed(MULT_83(18)(MULT_SIZE-1) & MULT_83(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(18)(MULT_SIZE-1) & MULT_84(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(19)<=signed(MULT_83(19)(MULT_SIZE-1) & MULT_83(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(19)(MULT_SIZE-1) & MULT_84(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(20)<=signed(MULT_83(20)(MULT_SIZE-1) & MULT_83(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(20)(MULT_SIZE-1) & MULT_84(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(21)<=signed(MULT_83(21)(MULT_SIZE-1) & MULT_83(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(21)(MULT_SIZE-1) & MULT_84(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(22)<=signed(MULT_83(22)(MULT_SIZE-1) & MULT_83(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(22)(MULT_SIZE-1) & MULT_84(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(23)<=signed(MULT_83(23)(MULT_SIZE-1) & MULT_83(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(23)(MULT_SIZE-1) & MULT_84(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(24)<=signed(MULT_83(24)(MULT_SIZE-1) & MULT_83(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(24)(MULT_SIZE-1) & MULT_84(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(25)<=signed(MULT_83(25)(MULT_SIZE-1) & MULT_83(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(25)(MULT_SIZE-1) & MULT_84(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(26)<=signed(MULT_83(26)(MULT_SIZE-1) & MULT_83(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(26)(MULT_SIZE-1) & MULT_84(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(27)<=signed(MULT_83(27)(MULT_SIZE-1) & MULT_83(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(27)(MULT_SIZE-1) & MULT_84(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(28)<=signed(MULT_83(28)(MULT_SIZE-1) & MULT_83(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(28)(MULT_SIZE-1) & MULT_84(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(29)<=signed(MULT_83(29)(MULT_SIZE-1) & MULT_83(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(29)(MULT_SIZE-1) & MULT_84(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(30)<=signed(MULT_83(30)(MULT_SIZE-1) & MULT_83(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(30)(MULT_SIZE-1) & MULT_84(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(31)<=signed(MULT_83(31)(MULT_SIZE-1) & MULT_83(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(31)(MULT_SIZE-1) & MULT_84(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(32)<=signed(MULT_83(32)(MULT_SIZE-1) & MULT_83(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(32)(MULT_SIZE-1) & MULT_84(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(33)<=signed(MULT_83(33)(MULT_SIZE-1) & MULT_83(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(33)(MULT_SIZE-1) & MULT_84(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(34)<=signed(MULT_83(34)(MULT_SIZE-1) & MULT_83(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(34)(MULT_SIZE-1) & MULT_84(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(35)<=signed(MULT_83(35)(MULT_SIZE-1) & MULT_83(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(35)(MULT_SIZE-1) & MULT_84(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(36)<=signed(MULT_83(36)(MULT_SIZE-1) & MULT_83(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(36)(MULT_SIZE-1) & MULT_84(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(37)<=signed(MULT_83(37)(MULT_SIZE-1) & MULT_83(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(37)(MULT_SIZE-1) & MULT_84(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(38)<=signed(MULT_83(38)(MULT_SIZE-1) & MULT_83(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(38)(MULT_SIZE-1) & MULT_84(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(39)<=signed(MULT_83(39)(MULT_SIZE-1) & MULT_83(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(39)(MULT_SIZE-1) & MULT_84(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(40)<=signed(MULT_83(40)(MULT_SIZE-1) & MULT_83(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(40)(MULT_SIZE-1) & MULT_84(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(41)<=signed(MULT_83(41)(MULT_SIZE-1) & MULT_83(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(41)(MULT_SIZE-1) & MULT_84(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(42)<=signed(MULT_83(42)(MULT_SIZE-1) & MULT_83(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(42)(MULT_SIZE-1) & MULT_84(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(43)<=signed(MULT_83(43)(MULT_SIZE-1) & MULT_83(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(43)(MULT_SIZE-1) & MULT_84(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(44)<=signed(MULT_83(44)(MULT_SIZE-1) & MULT_83(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(44)(MULT_SIZE-1) & MULT_84(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(45)<=signed(MULT_83(45)(MULT_SIZE-1) & MULT_83(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(45)(MULT_SIZE-1) & MULT_84(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(46)<=signed(MULT_83(46)(MULT_SIZE-1) & MULT_83(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(46)(MULT_SIZE-1) & MULT_84(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(47)<=signed(MULT_83(47)(MULT_SIZE-1) & MULT_83(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(47)(MULT_SIZE-1) & MULT_84(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(48)<=signed(MULT_83(48)(MULT_SIZE-1) & MULT_83(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(48)(MULT_SIZE-1) & MULT_84(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(49)<=signed(MULT_83(49)(MULT_SIZE-1) & MULT_83(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(49)(MULT_SIZE-1) & MULT_84(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(50)<=signed(MULT_83(50)(MULT_SIZE-1) & MULT_83(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(50)(MULT_SIZE-1) & MULT_84(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(51)<=signed(MULT_83(51)(MULT_SIZE-1) & MULT_83(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(51)(MULT_SIZE-1) & MULT_84(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(52)<=signed(MULT_83(52)(MULT_SIZE-1) & MULT_83(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(52)(MULT_SIZE-1) & MULT_84(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(53)<=signed(MULT_83(53)(MULT_SIZE-1) & MULT_83(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(53)(MULT_SIZE-1) & MULT_84(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(54)<=signed(MULT_83(54)(MULT_SIZE-1) & MULT_83(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(54)(MULT_SIZE-1) & MULT_84(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(55)<=signed(MULT_83(55)(MULT_SIZE-1) & MULT_83(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(55)(MULT_SIZE-1) & MULT_84(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(56)<=signed(MULT_83(56)(MULT_SIZE-1) & MULT_83(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(56)(MULT_SIZE-1) & MULT_84(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(57)<=signed(MULT_83(57)(MULT_SIZE-1) & MULT_83(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(57)(MULT_SIZE-1) & MULT_84(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(58)<=signed(MULT_83(58)(MULT_SIZE-1) & MULT_83(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(58)(MULT_SIZE-1) & MULT_84(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(59)<=signed(MULT_83(59)(MULT_SIZE-1) & MULT_83(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(59)(MULT_SIZE-1) & MULT_84(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(60)<=signed(MULT_83(60)(MULT_SIZE-1) & MULT_83(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(60)(MULT_SIZE-1) & MULT_84(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(61)<=signed(MULT_83(61)(MULT_SIZE-1) & MULT_83(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(61)(MULT_SIZE-1) & MULT_84(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(62)<=signed(MULT_83(62)(MULT_SIZE-1) & MULT_83(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(62)(MULT_SIZE-1) & MULT_84(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(63)<=signed(MULT_83(63)(MULT_SIZE-1) & MULT_83(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(63)(MULT_SIZE-1) & MULT_84(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(64)<=signed(MULT_83(64)(MULT_SIZE-1) & MULT_83(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(64)(MULT_SIZE-1) & MULT_84(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(65)<=signed(MULT_83(65)(MULT_SIZE-1) & MULT_83(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(65)(MULT_SIZE-1) & MULT_84(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(66)<=signed(MULT_83(66)(MULT_SIZE-1) & MULT_83(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(66)(MULT_SIZE-1) & MULT_84(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(67)<=signed(MULT_83(67)(MULT_SIZE-1) & MULT_83(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(67)(MULT_SIZE-1) & MULT_84(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(68)<=signed(MULT_83(68)(MULT_SIZE-1) & MULT_83(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(68)(MULT_SIZE-1) & MULT_84(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(69)<=signed(MULT_83(69)(MULT_SIZE-1) & MULT_83(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(69)(MULT_SIZE-1) & MULT_84(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(70)<=signed(MULT_83(70)(MULT_SIZE-1) & MULT_83(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(70)(MULT_SIZE-1) & MULT_84(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(71)<=signed(MULT_83(71)(MULT_SIZE-1) & MULT_83(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(71)(MULT_SIZE-1) & MULT_84(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(72)<=signed(MULT_83(72)(MULT_SIZE-1) & MULT_83(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(72)(MULT_SIZE-1) & MULT_84(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(73)<=signed(MULT_83(73)(MULT_SIZE-1) & MULT_83(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(73)(MULT_SIZE-1) & MULT_84(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(74)<=signed(MULT_83(74)(MULT_SIZE-1) & MULT_83(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(74)(MULT_SIZE-1) & MULT_84(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(75)<=signed(MULT_83(75)(MULT_SIZE-1) & MULT_83(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(75)(MULT_SIZE-1) & MULT_84(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(76)<=signed(MULT_83(76)(MULT_SIZE-1) & MULT_83(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(76)(MULT_SIZE-1) & MULT_84(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(77)<=signed(MULT_83(77)(MULT_SIZE-1) & MULT_83(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(77)(MULT_SIZE-1) & MULT_84(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(78)<=signed(MULT_83(78)(MULT_SIZE-1) & MULT_83(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(78)(MULT_SIZE-1) & MULT_84(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(79)<=signed(MULT_83(79)(MULT_SIZE-1) & MULT_83(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(79)(MULT_SIZE-1) & MULT_84(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(80)<=signed(MULT_83(80)(MULT_SIZE-1) & MULT_83(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(80)(MULT_SIZE-1) & MULT_84(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(81)<=signed(MULT_83(81)(MULT_SIZE-1) & MULT_83(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(81)(MULT_SIZE-1) & MULT_84(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(82)<=signed(MULT_83(82)(MULT_SIZE-1) & MULT_83(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(82)(MULT_SIZE-1) & MULT_84(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_42(83)<=signed(MULT_83(83)(MULT_SIZE-1) & MULT_83(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_84(83)(MULT_SIZE-1) & MULT_84(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_43(0)<=signed(MULT_85(0)(MULT_SIZE-1) & MULT_85(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(0)(MULT_SIZE-1) & MULT_86(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(1)<=signed(MULT_85(1)(MULT_SIZE-1) & MULT_85(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(1)(MULT_SIZE-1) & MULT_86(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(2)<=signed(MULT_85(2)(MULT_SIZE-1) & MULT_85(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(2)(MULT_SIZE-1) & MULT_86(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(3)<=signed(MULT_85(3)(MULT_SIZE-1) & MULT_85(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(3)(MULT_SIZE-1) & MULT_86(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(4)<=signed(MULT_85(4)(MULT_SIZE-1) & MULT_85(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(4)(MULT_SIZE-1) & MULT_86(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(5)<=signed(MULT_85(5)(MULT_SIZE-1) & MULT_85(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(5)(MULT_SIZE-1) & MULT_86(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(6)<=signed(MULT_85(6)(MULT_SIZE-1) & MULT_85(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(6)(MULT_SIZE-1) & MULT_86(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(7)<=signed(MULT_85(7)(MULT_SIZE-1) & MULT_85(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(7)(MULT_SIZE-1) & MULT_86(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(8)<=signed(MULT_85(8)(MULT_SIZE-1) & MULT_85(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(8)(MULT_SIZE-1) & MULT_86(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(9)<=signed(MULT_85(9)(MULT_SIZE-1) & MULT_85(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(9)(MULT_SIZE-1) & MULT_86(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(10)<=signed(MULT_85(10)(MULT_SIZE-1) & MULT_85(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(10)(MULT_SIZE-1) & MULT_86(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(11)<=signed(MULT_85(11)(MULT_SIZE-1) & MULT_85(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(11)(MULT_SIZE-1) & MULT_86(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(12)<=signed(MULT_85(12)(MULT_SIZE-1) & MULT_85(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(12)(MULT_SIZE-1) & MULT_86(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(13)<=signed(MULT_85(13)(MULT_SIZE-1) & MULT_85(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(13)(MULT_SIZE-1) & MULT_86(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(14)<=signed(MULT_85(14)(MULT_SIZE-1) & MULT_85(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(14)(MULT_SIZE-1) & MULT_86(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(15)<=signed(MULT_85(15)(MULT_SIZE-1) & MULT_85(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(15)(MULT_SIZE-1) & MULT_86(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(16)<=signed(MULT_85(16)(MULT_SIZE-1) & MULT_85(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(16)(MULT_SIZE-1) & MULT_86(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(17)<=signed(MULT_85(17)(MULT_SIZE-1) & MULT_85(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(17)(MULT_SIZE-1) & MULT_86(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(18)<=signed(MULT_85(18)(MULT_SIZE-1) & MULT_85(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(18)(MULT_SIZE-1) & MULT_86(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(19)<=signed(MULT_85(19)(MULT_SIZE-1) & MULT_85(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(19)(MULT_SIZE-1) & MULT_86(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(20)<=signed(MULT_85(20)(MULT_SIZE-1) & MULT_85(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(20)(MULT_SIZE-1) & MULT_86(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(21)<=signed(MULT_85(21)(MULT_SIZE-1) & MULT_85(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(21)(MULT_SIZE-1) & MULT_86(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(22)<=signed(MULT_85(22)(MULT_SIZE-1) & MULT_85(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(22)(MULT_SIZE-1) & MULT_86(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(23)<=signed(MULT_85(23)(MULT_SIZE-1) & MULT_85(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(23)(MULT_SIZE-1) & MULT_86(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(24)<=signed(MULT_85(24)(MULT_SIZE-1) & MULT_85(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(24)(MULT_SIZE-1) & MULT_86(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(25)<=signed(MULT_85(25)(MULT_SIZE-1) & MULT_85(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(25)(MULT_SIZE-1) & MULT_86(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(26)<=signed(MULT_85(26)(MULT_SIZE-1) & MULT_85(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(26)(MULT_SIZE-1) & MULT_86(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(27)<=signed(MULT_85(27)(MULT_SIZE-1) & MULT_85(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(27)(MULT_SIZE-1) & MULT_86(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(28)<=signed(MULT_85(28)(MULT_SIZE-1) & MULT_85(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(28)(MULT_SIZE-1) & MULT_86(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(29)<=signed(MULT_85(29)(MULT_SIZE-1) & MULT_85(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(29)(MULT_SIZE-1) & MULT_86(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(30)<=signed(MULT_85(30)(MULT_SIZE-1) & MULT_85(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(30)(MULT_SIZE-1) & MULT_86(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(31)<=signed(MULT_85(31)(MULT_SIZE-1) & MULT_85(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(31)(MULT_SIZE-1) & MULT_86(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(32)<=signed(MULT_85(32)(MULT_SIZE-1) & MULT_85(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(32)(MULT_SIZE-1) & MULT_86(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(33)<=signed(MULT_85(33)(MULT_SIZE-1) & MULT_85(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(33)(MULT_SIZE-1) & MULT_86(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(34)<=signed(MULT_85(34)(MULT_SIZE-1) & MULT_85(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(34)(MULT_SIZE-1) & MULT_86(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(35)<=signed(MULT_85(35)(MULT_SIZE-1) & MULT_85(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(35)(MULT_SIZE-1) & MULT_86(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(36)<=signed(MULT_85(36)(MULT_SIZE-1) & MULT_85(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(36)(MULT_SIZE-1) & MULT_86(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(37)<=signed(MULT_85(37)(MULT_SIZE-1) & MULT_85(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(37)(MULT_SIZE-1) & MULT_86(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(38)<=signed(MULT_85(38)(MULT_SIZE-1) & MULT_85(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(38)(MULT_SIZE-1) & MULT_86(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(39)<=signed(MULT_85(39)(MULT_SIZE-1) & MULT_85(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(39)(MULT_SIZE-1) & MULT_86(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(40)<=signed(MULT_85(40)(MULT_SIZE-1) & MULT_85(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(40)(MULT_SIZE-1) & MULT_86(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(41)<=signed(MULT_85(41)(MULT_SIZE-1) & MULT_85(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(41)(MULT_SIZE-1) & MULT_86(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(42)<=signed(MULT_85(42)(MULT_SIZE-1) & MULT_85(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(42)(MULT_SIZE-1) & MULT_86(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(43)<=signed(MULT_85(43)(MULT_SIZE-1) & MULT_85(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(43)(MULT_SIZE-1) & MULT_86(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(44)<=signed(MULT_85(44)(MULT_SIZE-1) & MULT_85(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(44)(MULT_SIZE-1) & MULT_86(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(45)<=signed(MULT_85(45)(MULT_SIZE-1) & MULT_85(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(45)(MULT_SIZE-1) & MULT_86(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(46)<=signed(MULT_85(46)(MULT_SIZE-1) & MULT_85(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(46)(MULT_SIZE-1) & MULT_86(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(47)<=signed(MULT_85(47)(MULT_SIZE-1) & MULT_85(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(47)(MULT_SIZE-1) & MULT_86(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(48)<=signed(MULT_85(48)(MULT_SIZE-1) & MULT_85(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(48)(MULT_SIZE-1) & MULT_86(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(49)<=signed(MULT_85(49)(MULT_SIZE-1) & MULT_85(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(49)(MULT_SIZE-1) & MULT_86(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(50)<=signed(MULT_85(50)(MULT_SIZE-1) & MULT_85(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(50)(MULT_SIZE-1) & MULT_86(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(51)<=signed(MULT_85(51)(MULT_SIZE-1) & MULT_85(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(51)(MULT_SIZE-1) & MULT_86(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(52)<=signed(MULT_85(52)(MULT_SIZE-1) & MULT_85(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(52)(MULT_SIZE-1) & MULT_86(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(53)<=signed(MULT_85(53)(MULT_SIZE-1) & MULT_85(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(53)(MULT_SIZE-1) & MULT_86(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(54)<=signed(MULT_85(54)(MULT_SIZE-1) & MULT_85(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(54)(MULT_SIZE-1) & MULT_86(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(55)<=signed(MULT_85(55)(MULT_SIZE-1) & MULT_85(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(55)(MULT_SIZE-1) & MULT_86(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(56)<=signed(MULT_85(56)(MULT_SIZE-1) & MULT_85(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(56)(MULT_SIZE-1) & MULT_86(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(57)<=signed(MULT_85(57)(MULT_SIZE-1) & MULT_85(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(57)(MULT_SIZE-1) & MULT_86(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(58)<=signed(MULT_85(58)(MULT_SIZE-1) & MULT_85(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(58)(MULT_SIZE-1) & MULT_86(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(59)<=signed(MULT_85(59)(MULT_SIZE-1) & MULT_85(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(59)(MULT_SIZE-1) & MULT_86(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(60)<=signed(MULT_85(60)(MULT_SIZE-1) & MULT_85(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(60)(MULT_SIZE-1) & MULT_86(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(61)<=signed(MULT_85(61)(MULT_SIZE-1) & MULT_85(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(61)(MULT_SIZE-1) & MULT_86(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(62)<=signed(MULT_85(62)(MULT_SIZE-1) & MULT_85(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(62)(MULT_SIZE-1) & MULT_86(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(63)<=signed(MULT_85(63)(MULT_SIZE-1) & MULT_85(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(63)(MULT_SIZE-1) & MULT_86(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(64)<=signed(MULT_85(64)(MULT_SIZE-1) & MULT_85(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(64)(MULT_SIZE-1) & MULT_86(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(65)<=signed(MULT_85(65)(MULT_SIZE-1) & MULT_85(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(65)(MULT_SIZE-1) & MULT_86(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(66)<=signed(MULT_85(66)(MULT_SIZE-1) & MULT_85(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(66)(MULT_SIZE-1) & MULT_86(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(67)<=signed(MULT_85(67)(MULT_SIZE-1) & MULT_85(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(67)(MULT_SIZE-1) & MULT_86(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(68)<=signed(MULT_85(68)(MULT_SIZE-1) & MULT_85(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(68)(MULT_SIZE-1) & MULT_86(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(69)<=signed(MULT_85(69)(MULT_SIZE-1) & MULT_85(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(69)(MULT_SIZE-1) & MULT_86(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(70)<=signed(MULT_85(70)(MULT_SIZE-1) & MULT_85(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(70)(MULT_SIZE-1) & MULT_86(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(71)<=signed(MULT_85(71)(MULT_SIZE-1) & MULT_85(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(71)(MULT_SIZE-1) & MULT_86(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(72)<=signed(MULT_85(72)(MULT_SIZE-1) & MULT_85(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(72)(MULT_SIZE-1) & MULT_86(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(73)<=signed(MULT_85(73)(MULT_SIZE-1) & MULT_85(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(73)(MULT_SIZE-1) & MULT_86(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(74)<=signed(MULT_85(74)(MULT_SIZE-1) & MULT_85(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(74)(MULT_SIZE-1) & MULT_86(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(75)<=signed(MULT_85(75)(MULT_SIZE-1) & MULT_85(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(75)(MULT_SIZE-1) & MULT_86(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(76)<=signed(MULT_85(76)(MULT_SIZE-1) & MULT_85(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(76)(MULT_SIZE-1) & MULT_86(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(77)<=signed(MULT_85(77)(MULT_SIZE-1) & MULT_85(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(77)(MULT_SIZE-1) & MULT_86(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(78)<=signed(MULT_85(78)(MULT_SIZE-1) & MULT_85(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(78)(MULT_SIZE-1) & MULT_86(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(79)<=signed(MULT_85(79)(MULT_SIZE-1) & MULT_85(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(79)(MULT_SIZE-1) & MULT_86(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(80)<=signed(MULT_85(80)(MULT_SIZE-1) & MULT_85(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(80)(MULT_SIZE-1) & MULT_86(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(81)<=signed(MULT_85(81)(MULT_SIZE-1) & MULT_85(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(81)(MULT_SIZE-1) & MULT_86(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(82)<=signed(MULT_85(82)(MULT_SIZE-1) & MULT_85(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(82)(MULT_SIZE-1) & MULT_86(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_43(83)<=signed(MULT_85(83)(MULT_SIZE-1) & MULT_85(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_86(83)(MULT_SIZE-1) & MULT_86(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_44(0)<=signed(MULT_87(0)(MULT_SIZE-1) & MULT_87(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(0)(MULT_SIZE-1) & MULT_88(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(1)<=signed(MULT_87(1)(MULT_SIZE-1) & MULT_87(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(1)(MULT_SIZE-1) & MULT_88(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(2)<=signed(MULT_87(2)(MULT_SIZE-1) & MULT_87(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(2)(MULT_SIZE-1) & MULT_88(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(3)<=signed(MULT_87(3)(MULT_SIZE-1) & MULT_87(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(3)(MULT_SIZE-1) & MULT_88(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(4)<=signed(MULT_87(4)(MULT_SIZE-1) & MULT_87(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(4)(MULT_SIZE-1) & MULT_88(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(5)<=signed(MULT_87(5)(MULT_SIZE-1) & MULT_87(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(5)(MULT_SIZE-1) & MULT_88(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(6)<=signed(MULT_87(6)(MULT_SIZE-1) & MULT_87(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(6)(MULT_SIZE-1) & MULT_88(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(7)<=signed(MULT_87(7)(MULT_SIZE-1) & MULT_87(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(7)(MULT_SIZE-1) & MULT_88(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(8)<=signed(MULT_87(8)(MULT_SIZE-1) & MULT_87(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(8)(MULT_SIZE-1) & MULT_88(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(9)<=signed(MULT_87(9)(MULT_SIZE-1) & MULT_87(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(9)(MULT_SIZE-1) & MULT_88(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(10)<=signed(MULT_87(10)(MULT_SIZE-1) & MULT_87(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(10)(MULT_SIZE-1) & MULT_88(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(11)<=signed(MULT_87(11)(MULT_SIZE-1) & MULT_87(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(11)(MULT_SIZE-1) & MULT_88(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(12)<=signed(MULT_87(12)(MULT_SIZE-1) & MULT_87(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(12)(MULT_SIZE-1) & MULT_88(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(13)<=signed(MULT_87(13)(MULT_SIZE-1) & MULT_87(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(13)(MULT_SIZE-1) & MULT_88(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(14)<=signed(MULT_87(14)(MULT_SIZE-1) & MULT_87(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(14)(MULT_SIZE-1) & MULT_88(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(15)<=signed(MULT_87(15)(MULT_SIZE-1) & MULT_87(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(15)(MULT_SIZE-1) & MULT_88(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(16)<=signed(MULT_87(16)(MULT_SIZE-1) & MULT_87(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(16)(MULT_SIZE-1) & MULT_88(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(17)<=signed(MULT_87(17)(MULT_SIZE-1) & MULT_87(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(17)(MULT_SIZE-1) & MULT_88(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(18)<=signed(MULT_87(18)(MULT_SIZE-1) & MULT_87(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(18)(MULT_SIZE-1) & MULT_88(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(19)<=signed(MULT_87(19)(MULT_SIZE-1) & MULT_87(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(19)(MULT_SIZE-1) & MULT_88(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(20)<=signed(MULT_87(20)(MULT_SIZE-1) & MULT_87(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(20)(MULT_SIZE-1) & MULT_88(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(21)<=signed(MULT_87(21)(MULT_SIZE-1) & MULT_87(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(21)(MULT_SIZE-1) & MULT_88(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(22)<=signed(MULT_87(22)(MULT_SIZE-1) & MULT_87(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(22)(MULT_SIZE-1) & MULT_88(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(23)<=signed(MULT_87(23)(MULT_SIZE-1) & MULT_87(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(23)(MULT_SIZE-1) & MULT_88(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(24)<=signed(MULT_87(24)(MULT_SIZE-1) & MULT_87(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(24)(MULT_SIZE-1) & MULT_88(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(25)<=signed(MULT_87(25)(MULT_SIZE-1) & MULT_87(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(25)(MULT_SIZE-1) & MULT_88(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(26)<=signed(MULT_87(26)(MULT_SIZE-1) & MULT_87(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(26)(MULT_SIZE-1) & MULT_88(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(27)<=signed(MULT_87(27)(MULT_SIZE-1) & MULT_87(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(27)(MULT_SIZE-1) & MULT_88(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(28)<=signed(MULT_87(28)(MULT_SIZE-1) & MULT_87(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(28)(MULT_SIZE-1) & MULT_88(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(29)<=signed(MULT_87(29)(MULT_SIZE-1) & MULT_87(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(29)(MULT_SIZE-1) & MULT_88(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(30)<=signed(MULT_87(30)(MULT_SIZE-1) & MULT_87(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(30)(MULT_SIZE-1) & MULT_88(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(31)<=signed(MULT_87(31)(MULT_SIZE-1) & MULT_87(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(31)(MULT_SIZE-1) & MULT_88(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(32)<=signed(MULT_87(32)(MULT_SIZE-1) & MULT_87(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(32)(MULT_SIZE-1) & MULT_88(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(33)<=signed(MULT_87(33)(MULT_SIZE-1) & MULT_87(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(33)(MULT_SIZE-1) & MULT_88(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(34)<=signed(MULT_87(34)(MULT_SIZE-1) & MULT_87(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(34)(MULT_SIZE-1) & MULT_88(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(35)<=signed(MULT_87(35)(MULT_SIZE-1) & MULT_87(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(35)(MULT_SIZE-1) & MULT_88(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(36)<=signed(MULT_87(36)(MULT_SIZE-1) & MULT_87(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(36)(MULT_SIZE-1) & MULT_88(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(37)<=signed(MULT_87(37)(MULT_SIZE-1) & MULT_87(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(37)(MULT_SIZE-1) & MULT_88(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(38)<=signed(MULT_87(38)(MULT_SIZE-1) & MULT_87(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(38)(MULT_SIZE-1) & MULT_88(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(39)<=signed(MULT_87(39)(MULT_SIZE-1) & MULT_87(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(39)(MULT_SIZE-1) & MULT_88(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(40)<=signed(MULT_87(40)(MULT_SIZE-1) & MULT_87(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(40)(MULT_SIZE-1) & MULT_88(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(41)<=signed(MULT_87(41)(MULT_SIZE-1) & MULT_87(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(41)(MULT_SIZE-1) & MULT_88(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(42)<=signed(MULT_87(42)(MULT_SIZE-1) & MULT_87(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(42)(MULT_SIZE-1) & MULT_88(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(43)<=signed(MULT_87(43)(MULT_SIZE-1) & MULT_87(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(43)(MULT_SIZE-1) & MULT_88(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(44)<=signed(MULT_87(44)(MULT_SIZE-1) & MULT_87(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(44)(MULT_SIZE-1) & MULT_88(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(45)<=signed(MULT_87(45)(MULT_SIZE-1) & MULT_87(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(45)(MULT_SIZE-1) & MULT_88(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(46)<=signed(MULT_87(46)(MULT_SIZE-1) & MULT_87(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(46)(MULT_SIZE-1) & MULT_88(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(47)<=signed(MULT_87(47)(MULT_SIZE-1) & MULT_87(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(47)(MULT_SIZE-1) & MULT_88(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(48)<=signed(MULT_87(48)(MULT_SIZE-1) & MULT_87(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(48)(MULT_SIZE-1) & MULT_88(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(49)<=signed(MULT_87(49)(MULT_SIZE-1) & MULT_87(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(49)(MULT_SIZE-1) & MULT_88(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(50)<=signed(MULT_87(50)(MULT_SIZE-1) & MULT_87(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(50)(MULT_SIZE-1) & MULT_88(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(51)<=signed(MULT_87(51)(MULT_SIZE-1) & MULT_87(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(51)(MULT_SIZE-1) & MULT_88(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(52)<=signed(MULT_87(52)(MULT_SIZE-1) & MULT_87(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(52)(MULT_SIZE-1) & MULT_88(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(53)<=signed(MULT_87(53)(MULT_SIZE-1) & MULT_87(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(53)(MULT_SIZE-1) & MULT_88(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(54)<=signed(MULT_87(54)(MULT_SIZE-1) & MULT_87(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(54)(MULT_SIZE-1) & MULT_88(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(55)<=signed(MULT_87(55)(MULT_SIZE-1) & MULT_87(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(55)(MULT_SIZE-1) & MULT_88(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(56)<=signed(MULT_87(56)(MULT_SIZE-1) & MULT_87(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(56)(MULT_SIZE-1) & MULT_88(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(57)<=signed(MULT_87(57)(MULT_SIZE-1) & MULT_87(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(57)(MULT_SIZE-1) & MULT_88(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(58)<=signed(MULT_87(58)(MULT_SIZE-1) & MULT_87(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(58)(MULT_SIZE-1) & MULT_88(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(59)<=signed(MULT_87(59)(MULT_SIZE-1) & MULT_87(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(59)(MULT_SIZE-1) & MULT_88(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(60)<=signed(MULT_87(60)(MULT_SIZE-1) & MULT_87(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(60)(MULT_SIZE-1) & MULT_88(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(61)<=signed(MULT_87(61)(MULT_SIZE-1) & MULT_87(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(61)(MULT_SIZE-1) & MULT_88(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(62)<=signed(MULT_87(62)(MULT_SIZE-1) & MULT_87(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(62)(MULT_SIZE-1) & MULT_88(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(63)<=signed(MULT_87(63)(MULT_SIZE-1) & MULT_87(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(63)(MULT_SIZE-1) & MULT_88(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(64)<=signed(MULT_87(64)(MULT_SIZE-1) & MULT_87(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(64)(MULT_SIZE-1) & MULT_88(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(65)<=signed(MULT_87(65)(MULT_SIZE-1) & MULT_87(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(65)(MULT_SIZE-1) & MULT_88(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(66)<=signed(MULT_87(66)(MULT_SIZE-1) & MULT_87(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(66)(MULT_SIZE-1) & MULT_88(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(67)<=signed(MULT_87(67)(MULT_SIZE-1) & MULT_87(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(67)(MULT_SIZE-1) & MULT_88(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(68)<=signed(MULT_87(68)(MULT_SIZE-1) & MULT_87(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(68)(MULT_SIZE-1) & MULT_88(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(69)<=signed(MULT_87(69)(MULT_SIZE-1) & MULT_87(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(69)(MULT_SIZE-1) & MULT_88(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(70)<=signed(MULT_87(70)(MULT_SIZE-1) & MULT_87(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(70)(MULT_SIZE-1) & MULT_88(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(71)<=signed(MULT_87(71)(MULT_SIZE-1) & MULT_87(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(71)(MULT_SIZE-1) & MULT_88(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(72)<=signed(MULT_87(72)(MULT_SIZE-1) & MULT_87(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(72)(MULT_SIZE-1) & MULT_88(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(73)<=signed(MULT_87(73)(MULT_SIZE-1) & MULT_87(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(73)(MULT_SIZE-1) & MULT_88(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(74)<=signed(MULT_87(74)(MULT_SIZE-1) & MULT_87(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(74)(MULT_SIZE-1) & MULT_88(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(75)<=signed(MULT_87(75)(MULT_SIZE-1) & MULT_87(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(75)(MULT_SIZE-1) & MULT_88(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(76)<=signed(MULT_87(76)(MULT_SIZE-1) & MULT_87(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(76)(MULT_SIZE-1) & MULT_88(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(77)<=signed(MULT_87(77)(MULT_SIZE-1) & MULT_87(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(77)(MULT_SIZE-1) & MULT_88(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(78)<=signed(MULT_87(78)(MULT_SIZE-1) & MULT_87(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(78)(MULT_SIZE-1) & MULT_88(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(79)<=signed(MULT_87(79)(MULT_SIZE-1) & MULT_87(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(79)(MULT_SIZE-1) & MULT_88(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(80)<=signed(MULT_87(80)(MULT_SIZE-1) & MULT_87(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(80)(MULT_SIZE-1) & MULT_88(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(81)<=signed(MULT_87(81)(MULT_SIZE-1) & MULT_87(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(81)(MULT_SIZE-1) & MULT_88(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(82)<=signed(MULT_87(82)(MULT_SIZE-1) & MULT_87(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(82)(MULT_SIZE-1) & MULT_88(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_44(83)<=signed(MULT_87(83)(MULT_SIZE-1) & MULT_87(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_88(83)(MULT_SIZE-1) & MULT_88(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_45(0)<=signed(MULT_89(0)(MULT_SIZE-1) & MULT_89(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(0)(MULT_SIZE-1) & MULT_90(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(1)<=signed(MULT_89(1)(MULT_SIZE-1) & MULT_89(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(1)(MULT_SIZE-1) & MULT_90(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(2)<=signed(MULT_89(2)(MULT_SIZE-1) & MULT_89(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(2)(MULT_SIZE-1) & MULT_90(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(3)<=signed(MULT_89(3)(MULT_SIZE-1) & MULT_89(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(3)(MULT_SIZE-1) & MULT_90(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(4)<=signed(MULT_89(4)(MULT_SIZE-1) & MULT_89(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(4)(MULT_SIZE-1) & MULT_90(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(5)<=signed(MULT_89(5)(MULT_SIZE-1) & MULT_89(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(5)(MULT_SIZE-1) & MULT_90(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(6)<=signed(MULT_89(6)(MULT_SIZE-1) & MULT_89(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(6)(MULT_SIZE-1) & MULT_90(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(7)<=signed(MULT_89(7)(MULT_SIZE-1) & MULT_89(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(7)(MULT_SIZE-1) & MULT_90(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(8)<=signed(MULT_89(8)(MULT_SIZE-1) & MULT_89(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(8)(MULT_SIZE-1) & MULT_90(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(9)<=signed(MULT_89(9)(MULT_SIZE-1) & MULT_89(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(9)(MULT_SIZE-1) & MULT_90(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(10)<=signed(MULT_89(10)(MULT_SIZE-1) & MULT_89(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(10)(MULT_SIZE-1) & MULT_90(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(11)<=signed(MULT_89(11)(MULT_SIZE-1) & MULT_89(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(11)(MULT_SIZE-1) & MULT_90(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(12)<=signed(MULT_89(12)(MULT_SIZE-1) & MULT_89(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(12)(MULT_SIZE-1) & MULT_90(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(13)<=signed(MULT_89(13)(MULT_SIZE-1) & MULT_89(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(13)(MULT_SIZE-1) & MULT_90(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(14)<=signed(MULT_89(14)(MULT_SIZE-1) & MULT_89(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(14)(MULT_SIZE-1) & MULT_90(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(15)<=signed(MULT_89(15)(MULT_SIZE-1) & MULT_89(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(15)(MULT_SIZE-1) & MULT_90(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(16)<=signed(MULT_89(16)(MULT_SIZE-1) & MULT_89(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(16)(MULT_SIZE-1) & MULT_90(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(17)<=signed(MULT_89(17)(MULT_SIZE-1) & MULT_89(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(17)(MULT_SIZE-1) & MULT_90(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(18)<=signed(MULT_89(18)(MULT_SIZE-1) & MULT_89(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(18)(MULT_SIZE-1) & MULT_90(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(19)<=signed(MULT_89(19)(MULT_SIZE-1) & MULT_89(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(19)(MULT_SIZE-1) & MULT_90(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(20)<=signed(MULT_89(20)(MULT_SIZE-1) & MULT_89(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(20)(MULT_SIZE-1) & MULT_90(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(21)<=signed(MULT_89(21)(MULT_SIZE-1) & MULT_89(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(21)(MULT_SIZE-1) & MULT_90(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(22)<=signed(MULT_89(22)(MULT_SIZE-1) & MULT_89(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(22)(MULT_SIZE-1) & MULT_90(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(23)<=signed(MULT_89(23)(MULT_SIZE-1) & MULT_89(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(23)(MULT_SIZE-1) & MULT_90(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(24)<=signed(MULT_89(24)(MULT_SIZE-1) & MULT_89(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(24)(MULT_SIZE-1) & MULT_90(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(25)<=signed(MULT_89(25)(MULT_SIZE-1) & MULT_89(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(25)(MULT_SIZE-1) & MULT_90(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(26)<=signed(MULT_89(26)(MULT_SIZE-1) & MULT_89(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(26)(MULT_SIZE-1) & MULT_90(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(27)<=signed(MULT_89(27)(MULT_SIZE-1) & MULT_89(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(27)(MULT_SIZE-1) & MULT_90(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(28)<=signed(MULT_89(28)(MULT_SIZE-1) & MULT_89(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(28)(MULT_SIZE-1) & MULT_90(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(29)<=signed(MULT_89(29)(MULT_SIZE-1) & MULT_89(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(29)(MULT_SIZE-1) & MULT_90(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(30)<=signed(MULT_89(30)(MULT_SIZE-1) & MULT_89(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(30)(MULT_SIZE-1) & MULT_90(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(31)<=signed(MULT_89(31)(MULT_SIZE-1) & MULT_89(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(31)(MULT_SIZE-1) & MULT_90(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(32)<=signed(MULT_89(32)(MULT_SIZE-1) & MULT_89(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(32)(MULT_SIZE-1) & MULT_90(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(33)<=signed(MULT_89(33)(MULT_SIZE-1) & MULT_89(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(33)(MULT_SIZE-1) & MULT_90(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(34)<=signed(MULT_89(34)(MULT_SIZE-1) & MULT_89(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(34)(MULT_SIZE-1) & MULT_90(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(35)<=signed(MULT_89(35)(MULT_SIZE-1) & MULT_89(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(35)(MULT_SIZE-1) & MULT_90(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(36)<=signed(MULT_89(36)(MULT_SIZE-1) & MULT_89(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(36)(MULT_SIZE-1) & MULT_90(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(37)<=signed(MULT_89(37)(MULT_SIZE-1) & MULT_89(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(37)(MULT_SIZE-1) & MULT_90(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(38)<=signed(MULT_89(38)(MULT_SIZE-1) & MULT_89(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(38)(MULT_SIZE-1) & MULT_90(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(39)<=signed(MULT_89(39)(MULT_SIZE-1) & MULT_89(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(39)(MULT_SIZE-1) & MULT_90(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(40)<=signed(MULT_89(40)(MULT_SIZE-1) & MULT_89(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(40)(MULT_SIZE-1) & MULT_90(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(41)<=signed(MULT_89(41)(MULT_SIZE-1) & MULT_89(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(41)(MULT_SIZE-1) & MULT_90(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(42)<=signed(MULT_89(42)(MULT_SIZE-1) & MULT_89(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(42)(MULT_SIZE-1) & MULT_90(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(43)<=signed(MULT_89(43)(MULT_SIZE-1) & MULT_89(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(43)(MULT_SIZE-1) & MULT_90(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(44)<=signed(MULT_89(44)(MULT_SIZE-1) & MULT_89(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(44)(MULT_SIZE-1) & MULT_90(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(45)<=signed(MULT_89(45)(MULT_SIZE-1) & MULT_89(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(45)(MULT_SIZE-1) & MULT_90(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(46)<=signed(MULT_89(46)(MULT_SIZE-1) & MULT_89(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(46)(MULT_SIZE-1) & MULT_90(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(47)<=signed(MULT_89(47)(MULT_SIZE-1) & MULT_89(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(47)(MULT_SIZE-1) & MULT_90(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(48)<=signed(MULT_89(48)(MULT_SIZE-1) & MULT_89(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(48)(MULT_SIZE-1) & MULT_90(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(49)<=signed(MULT_89(49)(MULT_SIZE-1) & MULT_89(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(49)(MULT_SIZE-1) & MULT_90(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(50)<=signed(MULT_89(50)(MULT_SIZE-1) & MULT_89(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(50)(MULT_SIZE-1) & MULT_90(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(51)<=signed(MULT_89(51)(MULT_SIZE-1) & MULT_89(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(51)(MULT_SIZE-1) & MULT_90(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(52)<=signed(MULT_89(52)(MULT_SIZE-1) & MULT_89(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(52)(MULT_SIZE-1) & MULT_90(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(53)<=signed(MULT_89(53)(MULT_SIZE-1) & MULT_89(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(53)(MULT_SIZE-1) & MULT_90(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(54)<=signed(MULT_89(54)(MULT_SIZE-1) & MULT_89(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(54)(MULT_SIZE-1) & MULT_90(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(55)<=signed(MULT_89(55)(MULT_SIZE-1) & MULT_89(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(55)(MULT_SIZE-1) & MULT_90(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(56)<=signed(MULT_89(56)(MULT_SIZE-1) & MULT_89(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(56)(MULT_SIZE-1) & MULT_90(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(57)<=signed(MULT_89(57)(MULT_SIZE-1) & MULT_89(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(57)(MULT_SIZE-1) & MULT_90(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(58)<=signed(MULT_89(58)(MULT_SIZE-1) & MULT_89(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(58)(MULT_SIZE-1) & MULT_90(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(59)<=signed(MULT_89(59)(MULT_SIZE-1) & MULT_89(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(59)(MULT_SIZE-1) & MULT_90(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(60)<=signed(MULT_89(60)(MULT_SIZE-1) & MULT_89(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(60)(MULT_SIZE-1) & MULT_90(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(61)<=signed(MULT_89(61)(MULT_SIZE-1) & MULT_89(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(61)(MULT_SIZE-1) & MULT_90(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(62)<=signed(MULT_89(62)(MULT_SIZE-1) & MULT_89(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(62)(MULT_SIZE-1) & MULT_90(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(63)<=signed(MULT_89(63)(MULT_SIZE-1) & MULT_89(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(63)(MULT_SIZE-1) & MULT_90(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(64)<=signed(MULT_89(64)(MULT_SIZE-1) & MULT_89(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(64)(MULT_SIZE-1) & MULT_90(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(65)<=signed(MULT_89(65)(MULT_SIZE-1) & MULT_89(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(65)(MULT_SIZE-1) & MULT_90(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(66)<=signed(MULT_89(66)(MULT_SIZE-1) & MULT_89(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(66)(MULT_SIZE-1) & MULT_90(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(67)<=signed(MULT_89(67)(MULT_SIZE-1) & MULT_89(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(67)(MULT_SIZE-1) & MULT_90(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(68)<=signed(MULT_89(68)(MULT_SIZE-1) & MULT_89(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(68)(MULT_SIZE-1) & MULT_90(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(69)<=signed(MULT_89(69)(MULT_SIZE-1) & MULT_89(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(69)(MULT_SIZE-1) & MULT_90(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(70)<=signed(MULT_89(70)(MULT_SIZE-1) & MULT_89(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(70)(MULT_SIZE-1) & MULT_90(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(71)<=signed(MULT_89(71)(MULT_SIZE-1) & MULT_89(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(71)(MULT_SIZE-1) & MULT_90(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(72)<=signed(MULT_89(72)(MULT_SIZE-1) & MULT_89(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(72)(MULT_SIZE-1) & MULT_90(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(73)<=signed(MULT_89(73)(MULT_SIZE-1) & MULT_89(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(73)(MULT_SIZE-1) & MULT_90(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(74)<=signed(MULT_89(74)(MULT_SIZE-1) & MULT_89(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(74)(MULT_SIZE-1) & MULT_90(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(75)<=signed(MULT_89(75)(MULT_SIZE-1) & MULT_89(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(75)(MULT_SIZE-1) & MULT_90(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(76)<=signed(MULT_89(76)(MULT_SIZE-1) & MULT_89(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(76)(MULT_SIZE-1) & MULT_90(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(77)<=signed(MULT_89(77)(MULT_SIZE-1) & MULT_89(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(77)(MULT_SIZE-1) & MULT_90(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(78)<=signed(MULT_89(78)(MULT_SIZE-1) & MULT_89(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(78)(MULT_SIZE-1) & MULT_90(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(79)<=signed(MULT_89(79)(MULT_SIZE-1) & MULT_89(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(79)(MULT_SIZE-1) & MULT_90(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(80)<=signed(MULT_89(80)(MULT_SIZE-1) & MULT_89(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(80)(MULT_SIZE-1) & MULT_90(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(81)<=signed(MULT_89(81)(MULT_SIZE-1) & MULT_89(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(81)(MULT_SIZE-1) & MULT_90(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(82)<=signed(MULT_89(82)(MULT_SIZE-1) & MULT_89(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(82)(MULT_SIZE-1) & MULT_90(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_45(83)<=signed(MULT_89(83)(MULT_SIZE-1) & MULT_89(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_90(83)(MULT_SIZE-1) & MULT_90(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_46(0)<=signed(MULT_91(0)(MULT_SIZE-1) & MULT_91(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(0)(MULT_SIZE-1) & MULT_92(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(1)<=signed(MULT_91(1)(MULT_SIZE-1) & MULT_91(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(1)(MULT_SIZE-1) & MULT_92(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(2)<=signed(MULT_91(2)(MULT_SIZE-1) & MULT_91(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(2)(MULT_SIZE-1) & MULT_92(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(3)<=signed(MULT_91(3)(MULT_SIZE-1) & MULT_91(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(3)(MULT_SIZE-1) & MULT_92(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(4)<=signed(MULT_91(4)(MULT_SIZE-1) & MULT_91(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(4)(MULT_SIZE-1) & MULT_92(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(5)<=signed(MULT_91(5)(MULT_SIZE-1) & MULT_91(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(5)(MULT_SIZE-1) & MULT_92(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(6)<=signed(MULT_91(6)(MULT_SIZE-1) & MULT_91(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(6)(MULT_SIZE-1) & MULT_92(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(7)<=signed(MULT_91(7)(MULT_SIZE-1) & MULT_91(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(7)(MULT_SIZE-1) & MULT_92(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(8)<=signed(MULT_91(8)(MULT_SIZE-1) & MULT_91(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(8)(MULT_SIZE-1) & MULT_92(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(9)<=signed(MULT_91(9)(MULT_SIZE-1) & MULT_91(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(9)(MULT_SIZE-1) & MULT_92(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(10)<=signed(MULT_91(10)(MULT_SIZE-1) & MULT_91(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(10)(MULT_SIZE-1) & MULT_92(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(11)<=signed(MULT_91(11)(MULT_SIZE-1) & MULT_91(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(11)(MULT_SIZE-1) & MULT_92(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(12)<=signed(MULT_91(12)(MULT_SIZE-1) & MULT_91(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(12)(MULT_SIZE-1) & MULT_92(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(13)<=signed(MULT_91(13)(MULT_SIZE-1) & MULT_91(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(13)(MULT_SIZE-1) & MULT_92(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(14)<=signed(MULT_91(14)(MULT_SIZE-1) & MULT_91(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(14)(MULT_SIZE-1) & MULT_92(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(15)<=signed(MULT_91(15)(MULT_SIZE-1) & MULT_91(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(15)(MULT_SIZE-1) & MULT_92(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(16)<=signed(MULT_91(16)(MULT_SIZE-1) & MULT_91(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(16)(MULT_SIZE-1) & MULT_92(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(17)<=signed(MULT_91(17)(MULT_SIZE-1) & MULT_91(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(17)(MULT_SIZE-1) & MULT_92(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(18)<=signed(MULT_91(18)(MULT_SIZE-1) & MULT_91(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(18)(MULT_SIZE-1) & MULT_92(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(19)<=signed(MULT_91(19)(MULT_SIZE-1) & MULT_91(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(19)(MULT_SIZE-1) & MULT_92(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(20)<=signed(MULT_91(20)(MULT_SIZE-1) & MULT_91(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(20)(MULT_SIZE-1) & MULT_92(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(21)<=signed(MULT_91(21)(MULT_SIZE-1) & MULT_91(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(21)(MULT_SIZE-1) & MULT_92(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(22)<=signed(MULT_91(22)(MULT_SIZE-1) & MULT_91(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(22)(MULT_SIZE-1) & MULT_92(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(23)<=signed(MULT_91(23)(MULT_SIZE-1) & MULT_91(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(23)(MULT_SIZE-1) & MULT_92(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(24)<=signed(MULT_91(24)(MULT_SIZE-1) & MULT_91(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(24)(MULT_SIZE-1) & MULT_92(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(25)<=signed(MULT_91(25)(MULT_SIZE-1) & MULT_91(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(25)(MULT_SIZE-1) & MULT_92(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(26)<=signed(MULT_91(26)(MULT_SIZE-1) & MULT_91(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(26)(MULT_SIZE-1) & MULT_92(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(27)<=signed(MULT_91(27)(MULT_SIZE-1) & MULT_91(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(27)(MULT_SIZE-1) & MULT_92(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(28)<=signed(MULT_91(28)(MULT_SIZE-1) & MULT_91(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(28)(MULT_SIZE-1) & MULT_92(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(29)<=signed(MULT_91(29)(MULT_SIZE-1) & MULT_91(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(29)(MULT_SIZE-1) & MULT_92(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(30)<=signed(MULT_91(30)(MULT_SIZE-1) & MULT_91(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(30)(MULT_SIZE-1) & MULT_92(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(31)<=signed(MULT_91(31)(MULT_SIZE-1) & MULT_91(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(31)(MULT_SIZE-1) & MULT_92(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(32)<=signed(MULT_91(32)(MULT_SIZE-1) & MULT_91(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(32)(MULT_SIZE-1) & MULT_92(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(33)<=signed(MULT_91(33)(MULT_SIZE-1) & MULT_91(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(33)(MULT_SIZE-1) & MULT_92(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(34)<=signed(MULT_91(34)(MULT_SIZE-1) & MULT_91(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(34)(MULT_SIZE-1) & MULT_92(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(35)<=signed(MULT_91(35)(MULT_SIZE-1) & MULT_91(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(35)(MULT_SIZE-1) & MULT_92(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(36)<=signed(MULT_91(36)(MULT_SIZE-1) & MULT_91(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(36)(MULT_SIZE-1) & MULT_92(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(37)<=signed(MULT_91(37)(MULT_SIZE-1) & MULT_91(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(37)(MULT_SIZE-1) & MULT_92(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(38)<=signed(MULT_91(38)(MULT_SIZE-1) & MULT_91(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(38)(MULT_SIZE-1) & MULT_92(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(39)<=signed(MULT_91(39)(MULT_SIZE-1) & MULT_91(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(39)(MULT_SIZE-1) & MULT_92(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(40)<=signed(MULT_91(40)(MULT_SIZE-1) & MULT_91(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(40)(MULT_SIZE-1) & MULT_92(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(41)<=signed(MULT_91(41)(MULT_SIZE-1) & MULT_91(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(41)(MULT_SIZE-1) & MULT_92(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(42)<=signed(MULT_91(42)(MULT_SIZE-1) & MULT_91(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(42)(MULT_SIZE-1) & MULT_92(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(43)<=signed(MULT_91(43)(MULT_SIZE-1) & MULT_91(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(43)(MULT_SIZE-1) & MULT_92(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(44)<=signed(MULT_91(44)(MULT_SIZE-1) & MULT_91(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(44)(MULT_SIZE-1) & MULT_92(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(45)<=signed(MULT_91(45)(MULT_SIZE-1) & MULT_91(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(45)(MULT_SIZE-1) & MULT_92(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(46)<=signed(MULT_91(46)(MULT_SIZE-1) & MULT_91(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(46)(MULT_SIZE-1) & MULT_92(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(47)<=signed(MULT_91(47)(MULT_SIZE-1) & MULT_91(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(47)(MULT_SIZE-1) & MULT_92(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(48)<=signed(MULT_91(48)(MULT_SIZE-1) & MULT_91(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(48)(MULT_SIZE-1) & MULT_92(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(49)<=signed(MULT_91(49)(MULT_SIZE-1) & MULT_91(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(49)(MULT_SIZE-1) & MULT_92(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(50)<=signed(MULT_91(50)(MULT_SIZE-1) & MULT_91(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(50)(MULT_SIZE-1) & MULT_92(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(51)<=signed(MULT_91(51)(MULT_SIZE-1) & MULT_91(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(51)(MULT_SIZE-1) & MULT_92(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(52)<=signed(MULT_91(52)(MULT_SIZE-1) & MULT_91(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(52)(MULT_SIZE-1) & MULT_92(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(53)<=signed(MULT_91(53)(MULT_SIZE-1) & MULT_91(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(53)(MULT_SIZE-1) & MULT_92(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(54)<=signed(MULT_91(54)(MULT_SIZE-1) & MULT_91(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(54)(MULT_SIZE-1) & MULT_92(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(55)<=signed(MULT_91(55)(MULT_SIZE-1) & MULT_91(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(55)(MULT_SIZE-1) & MULT_92(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(56)<=signed(MULT_91(56)(MULT_SIZE-1) & MULT_91(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(56)(MULT_SIZE-1) & MULT_92(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(57)<=signed(MULT_91(57)(MULT_SIZE-1) & MULT_91(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(57)(MULT_SIZE-1) & MULT_92(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(58)<=signed(MULT_91(58)(MULT_SIZE-1) & MULT_91(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(58)(MULT_SIZE-1) & MULT_92(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(59)<=signed(MULT_91(59)(MULT_SIZE-1) & MULT_91(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(59)(MULT_SIZE-1) & MULT_92(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(60)<=signed(MULT_91(60)(MULT_SIZE-1) & MULT_91(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(60)(MULT_SIZE-1) & MULT_92(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(61)<=signed(MULT_91(61)(MULT_SIZE-1) & MULT_91(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(61)(MULT_SIZE-1) & MULT_92(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(62)<=signed(MULT_91(62)(MULT_SIZE-1) & MULT_91(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(62)(MULT_SIZE-1) & MULT_92(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(63)<=signed(MULT_91(63)(MULT_SIZE-1) & MULT_91(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(63)(MULT_SIZE-1) & MULT_92(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(64)<=signed(MULT_91(64)(MULT_SIZE-1) & MULT_91(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(64)(MULT_SIZE-1) & MULT_92(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(65)<=signed(MULT_91(65)(MULT_SIZE-1) & MULT_91(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(65)(MULT_SIZE-1) & MULT_92(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(66)<=signed(MULT_91(66)(MULT_SIZE-1) & MULT_91(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(66)(MULT_SIZE-1) & MULT_92(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(67)<=signed(MULT_91(67)(MULT_SIZE-1) & MULT_91(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(67)(MULT_SIZE-1) & MULT_92(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(68)<=signed(MULT_91(68)(MULT_SIZE-1) & MULT_91(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(68)(MULT_SIZE-1) & MULT_92(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(69)<=signed(MULT_91(69)(MULT_SIZE-1) & MULT_91(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(69)(MULT_SIZE-1) & MULT_92(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(70)<=signed(MULT_91(70)(MULT_SIZE-1) & MULT_91(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(70)(MULT_SIZE-1) & MULT_92(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(71)<=signed(MULT_91(71)(MULT_SIZE-1) & MULT_91(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(71)(MULT_SIZE-1) & MULT_92(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(72)<=signed(MULT_91(72)(MULT_SIZE-1) & MULT_91(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(72)(MULT_SIZE-1) & MULT_92(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(73)<=signed(MULT_91(73)(MULT_SIZE-1) & MULT_91(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(73)(MULT_SIZE-1) & MULT_92(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(74)<=signed(MULT_91(74)(MULT_SIZE-1) & MULT_91(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(74)(MULT_SIZE-1) & MULT_92(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(75)<=signed(MULT_91(75)(MULT_SIZE-1) & MULT_91(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(75)(MULT_SIZE-1) & MULT_92(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(76)<=signed(MULT_91(76)(MULT_SIZE-1) & MULT_91(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(76)(MULT_SIZE-1) & MULT_92(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(77)<=signed(MULT_91(77)(MULT_SIZE-1) & MULT_91(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(77)(MULT_SIZE-1) & MULT_92(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(78)<=signed(MULT_91(78)(MULT_SIZE-1) & MULT_91(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(78)(MULT_SIZE-1) & MULT_92(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(79)<=signed(MULT_91(79)(MULT_SIZE-1) & MULT_91(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(79)(MULT_SIZE-1) & MULT_92(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(80)<=signed(MULT_91(80)(MULT_SIZE-1) & MULT_91(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(80)(MULT_SIZE-1) & MULT_92(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(81)<=signed(MULT_91(81)(MULT_SIZE-1) & MULT_91(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(81)(MULT_SIZE-1) & MULT_92(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(82)<=signed(MULT_91(82)(MULT_SIZE-1) & MULT_91(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(82)(MULT_SIZE-1) & MULT_92(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_46(83)<=signed(MULT_91(83)(MULT_SIZE-1) & MULT_91(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_92(83)(MULT_SIZE-1) & MULT_92(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_47(0)<=signed(MULT_93(0)(MULT_SIZE-1) & MULT_93(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(0)(MULT_SIZE-1) & MULT_94(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(1)<=signed(MULT_93(1)(MULT_SIZE-1) & MULT_93(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(1)(MULT_SIZE-1) & MULT_94(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(2)<=signed(MULT_93(2)(MULT_SIZE-1) & MULT_93(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(2)(MULT_SIZE-1) & MULT_94(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(3)<=signed(MULT_93(3)(MULT_SIZE-1) & MULT_93(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(3)(MULT_SIZE-1) & MULT_94(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(4)<=signed(MULT_93(4)(MULT_SIZE-1) & MULT_93(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(4)(MULT_SIZE-1) & MULT_94(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(5)<=signed(MULT_93(5)(MULT_SIZE-1) & MULT_93(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(5)(MULT_SIZE-1) & MULT_94(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(6)<=signed(MULT_93(6)(MULT_SIZE-1) & MULT_93(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(6)(MULT_SIZE-1) & MULT_94(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(7)<=signed(MULT_93(7)(MULT_SIZE-1) & MULT_93(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(7)(MULT_SIZE-1) & MULT_94(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(8)<=signed(MULT_93(8)(MULT_SIZE-1) & MULT_93(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(8)(MULT_SIZE-1) & MULT_94(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(9)<=signed(MULT_93(9)(MULT_SIZE-1) & MULT_93(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(9)(MULT_SIZE-1) & MULT_94(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(10)<=signed(MULT_93(10)(MULT_SIZE-1) & MULT_93(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(10)(MULT_SIZE-1) & MULT_94(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(11)<=signed(MULT_93(11)(MULT_SIZE-1) & MULT_93(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(11)(MULT_SIZE-1) & MULT_94(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(12)<=signed(MULT_93(12)(MULT_SIZE-1) & MULT_93(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(12)(MULT_SIZE-1) & MULT_94(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(13)<=signed(MULT_93(13)(MULT_SIZE-1) & MULT_93(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(13)(MULT_SIZE-1) & MULT_94(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(14)<=signed(MULT_93(14)(MULT_SIZE-1) & MULT_93(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(14)(MULT_SIZE-1) & MULT_94(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(15)<=signed(MULT_93(15)(MULT_SIZE-1) & MULT_93(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(15)(MULT_SIZE-1) & MULT_94(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(16)<=signed(MULT_93(16)(MULT_SIZE-1) & MULT_93(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(16)(MULT_SIZE-1) & MULT_94(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(17)<=signed(MULT_93(17)(MULT_SIZE-1) & MULT_93(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(17)(MULT_SIZE-1) & MULT_94(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(18)<=signed(MULT_93(18)(MULT_SIZE-1) & MULT_93(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(18)(MULT_SIZE-1) & MULT_94(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(19)<=signed(MULT_93(19)(MULT_SIZE-1) & MULT_93(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(19)(MULT_SIZE-1) & MULT_94(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(20)<=signed(MULT_93(20)(MULT_SIZE-1) & MULT_93(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(20)(MULT_SIZE-1) & MULT_94(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(21)<=signed(MULT_93(21)(MULT_SIZE-1) & MULT_93(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(21)(MULT_SIZE-1) & MULT_94(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(22)<=signed(MULT_93(22)(MULT_SIZE-1) & MULT_93(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(22)(MULT_SIZE-1) & MULT_94(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(23)<=signed(MULT_93(23)(MULT_SIZE-1) & MULT_93(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(23)(MULT_SIZE-1) & MULT_94(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(24)<=signed(MULT_93(24)(MULT_SIZE-1) & MULT_93(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(24)(MULT_SIZE-1) & MULT_94(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(25)<=signed(MULT_93(25)(MULT_SIZE-1) & MULT_93(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(25)(MULT_SIZE-1) & MULT_94(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(26)<=signed(MULT_93(26)(MULT_SIZE-1) & MULT_93(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(26)(MULT_SIZE-1) & MULT_94(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(27)<=signed(MULT_93(27)(MULT_SIZE-1) & MULT_93(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(27)(MULT_SIZE-1) & MULT_94(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(28)<=signed(MULT_93(28)(MULT_SIZE-1) & MULT_93(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(28)(MULT_SIZE-1) & MULT_94(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(29)<=signed(MULT_93(29)(MULT_SIZE-1) & MULT_93(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(29)(MULT_SIZE-1) & MULT_94(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(30)<=signed(MULT_93(30)(MULT_SIZE-1) & MULT_93(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(30)(MULT_SIZE-1) & MULT_94(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(31)<=signed(MULT_93(31)(MULT_SIZE-1) & MULT_93(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(31)(MULT_SIZE-1) & MULT_94(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(32)<=signed(MULT_93(32)(MULT_SIZE-1) & MULT_93(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(32)(MULT_SIZE-1) & MULT_94(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(33)<=signed(MULT_93(33)(MULT_SIZE-1) & MULT_93(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(33)(MULT_SIZE-1) & MULT_94(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(34)<=signed(MULT_93(34)(MULT_SIZE-1) & MULT_93(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(34)(MULT_SIZE-1) & MULT_94(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(35)<=signed(MULT_93(35)(MULT_SIZE-1) & MULT_93(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(35)(MULT_SIZE-1) & MULT_94(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(36)<=signed(MULT_93(36)(MULT_SIZE-1) & MULT_93(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(36)(MULT_SIZE-1) & MULT_94(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(37)<=signed(MULT_93(37)(MULT_SIZE-1) & MULT_93(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(37)(MULT_SIZE-1) & MULT_94(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(38)<=signed(MULT_93(38)(MULT_SIZE-1) & MULT_93(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(38)(MULT_SIZE-1) & MULT_94(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(39)<=signed(MULT_93(39)(MULT_SIZE-1) & MULT_93(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(39)(MULT_SIZE-1) & MULT_94(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(40)<=signed(MULT_93(40)(MULT_SIZE-1) & MULT_93(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(40)(MULT_SIZE-1) & MULT_94(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(41)<=signed(MULT_93(41)(MULT_SIZE-1) & MULT_93(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(41)(MULT_SIZE-1) & MULT_94(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(42)<=signed(MULT_93(42)(MULT_SIZE-1) & MULT_93(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(42)(MULT_SIZE-1) & MULT_94(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(43)<=signed(MULT_93(43)(MULT_SIZE-1) & MULT_93(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(43)(MULT_SIZE-1) & MULT_94(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(44)<=signed(MULT_93(44)(MULT_SIZE-1) & MULT_93(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(44)(MULT_SIZE-1) & MULT_94(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(45)<=signed(MULT_93(45)(MULT_SIZE-1) & MULT_93(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(45)(MULT_SIZE-1) & MULT_94(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(46)<=signed(MULT_93(46)(MULT_SIZE-1) & MULT_93(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(46)(MULT_SIZE-1) & MULT_94(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(47)<=signed(MULT_93(47)(MULT_SIZE-1) & MULT_93(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(47)(MULT_SIZE-1) & MULT_94(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(48)<=signed(MULT_93(48)(MULT_SIZE-1) & MULT_93(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(48)(MULT_SIZE-1) & MULT_94(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(49)<=signed(MULT_93(49)(MULT_SIZE-1) & MULT_93(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(49)(MULT_SIZE-1) & MULT_94(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(50)<=signed(MULT_93(50)(MULT_SIZE-1) & MULT_93(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(50)(MULT_SIZE-1) & MULT_94(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(51)<=signed(MULT_93(51)(MULT_SIZE-1) & MULT_93(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(51)(MULT_SIZE-1) & MULT_94(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(52)<=signed(MULT_93(52)(MULT_SIZE-1) & MULT_93(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(52)(MULT_SIZE-1) & MULT_94(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(53)<=signed(MULT_93(53)(MULT_SIZE-1) & MULT_93(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(53)(MULT_SIZE-1) & MULT_94(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(54)<=signed(MULT_93(54)(MULT_SIZE-1) & MULT_93(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(54)(MULT_SIZE-1) & MULT_94(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(55)<=signed(MULT_93(55)(MULT_SIZE-1) & MULT_93(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(55)(MULT_SIZE-1) & MULT_94(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(56)<=signed(MULT_93(56)(MULT_SIZE-1) & MULT_93(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(56)(MULT_SIZE-1) & MULT_94(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(57)<=signed(MULT_93(57)(MULT_SIZE-1) & MULT_93(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(57)(MULT_SIZE-1) & MULT_94(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(58)<=signed(MULT_93(58)(MULT_SIZE-1) & MULT_93(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(58)(MULT_SIZE-1) & MULT_94(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(59)<=signed(MULT_93(59)(MULT_SIZE-1) & MULT_93(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(59)(MULT_SIZE-1) & MULT_94(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(60)<=signed(MULT_93(60)(MULT_SIZE-1) & MULT_93(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(60)(MULT_SIZE-1) & MULT_94(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(61)<=signed(MULT_93(61)(MULT_SIZE-1) & MULT_93(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(61)(MULT_SIZE-1) & MULT_94(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(62)<=signed(MULT_93(62)(MULT_SIZE-1) & MULT_93(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(62)(MULT_SIZE-1) & MULT_94(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(63)<=signed(MULT_93(63)(MULT_SIZE-1) & MULT_93(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(63)(MULT_SIZE-1) & MULT_94(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(64)<=signed(MULT_93(64)(MULT_SIZE-1) & MULT_93(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(64)(MULT_SIZE-1) & MULT_94(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(65)<=signed(MULT_93(65)(MULT_SIZE-1) & MULT_93(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(65)(MULT_SIZE-1) & MULT_94(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(66)<=signed(MULT_93(66)(MULT_SIZE-1) & MULT_93(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(66)(MULT_SIZE-1) & MULT_94(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(67)<=signed(MULT_93(67)(MULT_SIZE-1) & MULT_93(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(67)(MULT_SIZE-1) & MULT_94(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(68)<=signed(MULT_93(68)(MULT_SIZE-1) & MULT_93(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(68)(MULT_SIZE-1) & MULT_94(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(69)<=signed(MULT_93(69)(MULT_SIZE-1) & MULT_93(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(69)(MULT_SIZE-1) & MULT_94(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(70)<=signed(MULT_93(70)(MULT_SIZE-1) & MULT_93(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(70)(MULT_SIZE-1) & MULT_94(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(71)<=signed(MULT_93(71)(MULT_SIZE-1) & MULT_93(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(71)(MULT_SIZE-1) & MULT_94(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(72)<=signed(MULT_93(72)(MULT_SIZE-1) & MULT_93(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(72)(MULT_SIZE-1) & MULT_94(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(73)<=signed(MULT_93(73)(MULT_SIZE-1) & MULT_93(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(73)(MULT_SIZE-1) & MULT_94(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(74)<=signed(MULT_93(74)(MULT_SIZE-1) & MULT_93(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(74)(MULT_SIZE-1) & MULT_94(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(75)<=signed(MULT_93(75)(MULT_SIZE-1) & MULT_93(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(75)(MULT_SIZE-1) & MULT_94(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(76)<=signed(MULT_93(76)(MULT_SIZE-1) & MULT_93(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(76)(MULT_SIZE-1) & MULT_94(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(77)<=signed(MULT_93(77)(MULT_SIZE-1) & MULT_93(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(77)(MULT_SIZE-1) & MULT_94(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(78)<=signed(MULT_93(78)(MULT_SIZE-1) & MULT_93(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(78)(MULT_SIZE-1) & MULT_94(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(79)<=signed(MULT_93(79)(MULT_SIZE-1) & MULT_93(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(79)(MULT_SIZE-1) & MULT_94(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(80)<=signed(MULT_93(80)(MULT_SIZE-1) & MULT_93(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(80)(MULT_SIZE-1) & MULT_94(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(81)<=signed(MULT_93(81)(MULT_SIZE-1) & MULT_93(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(81)(MULT_SIZE-1) & MULT_94(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(82)<=signed(MULT_93(82)(MULT_SIZE-1) & MULT_93(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(82)(MULT_SIZE-1) & MULT_94(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_47(83)<=signed(MULT_93(83)(MULT_SIZE-1) & MULT_93(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_94(83)(MULT_SIZE-1) & MULT_94(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_48(0)<=signed(MULT_95(0)(MULT_SIZE-1) & MULT_95(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(0)(MULT_SIZE-1) & MULT_96(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(1)<=signed(MULT_95(1)(MULT_SIZE-1) & MULT_95(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(1)(MULT_SIZE-1) & MULT_96(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(2)<=signed(MULT_95(2)(MULT_SIZE-1) & MULT_95(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(2)(MULT_SIZE-1) & MULT_96(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(3)<=signed(MULT_95(3)(MULT_SIZE-1) & MULT_95(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(3)(MULT_SIZE-1) & MULT_96(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(4)<=signed(MULT_95(4)(MULT_SIZE-1) & MULT_95(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(4)(MULT_SIZE-1) & MULT_96(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(5)<=signed(MULT_95(5)(MULT_SIZE-1) & MULT_95(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(5)(MULT_SIZE-1) & MULT_96(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(6)<=signed(MULT_95(6)(MULT_SIZE-1) & MULT_95(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(6)(MULT_SIZE-1) & MULT_96(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(7)<=signed(MULT_95(7)(MULT_SIZE-1) & MULT_95(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(7)(MULT_SIZE-1) & MULT_96(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(8)<=signed(MULT_95(8)(MULT_SIZE-1) & MULT_95(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(8)(MULT_SIZE-1) & MULT_96(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(9)<=signed(MULT_95(9)(MULT_SIZE-1) & MULT_95(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(9)(MULT_SIZE-1) & MULT_96(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(10)<=signed(MULT_95(10)(MULT_SIZE-1) & MULT_95(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(10)(MULT_SIZE-1) & MULT_96(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(11)<=signed(MULT_95(11)(MULT_SIZE-1) & MULT_95(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(11)(MULT_SIZE-1) & MULT_96(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(12)<=signed(MULT_95(12)(MULT_SIZE-1) & MULT_95(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(12)(MULT_SIZE-1) & MULT_96(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(13)<=signed(MULT_95(13)(MULT_SIZE-1) & MULT_95(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(13)(MULT_SIZE-1) & MULT_96(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(14)<=signed(MULT_95(14)(MULT_SIZE-1) & MULT_95(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(14)(MULT_SIZE-1) & MULT_96(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(15)<=signed(MULT_95(15)(MULT_SIZE-1) & MULT_95(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(15)(MULT_SIZE-1) & MULT_96(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(16)<=signed(MULT_95(16)(MULT_SIZE-1) & MULT_95(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(16)(MULT_SIZE-1) & MULT_96(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(17)<=signed(MULT_95(17)(MULT_SIZE-1) & MULT_95(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(17)(MULT_SIZE-1) & MULT_96(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(18)<=signed(MULT_95(18)(MULT_SIZE-1) & MULT_95(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(18)(MULT_SIZE-1) & MULT_96(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(19)<=signed(MULT_95(19)(MULT_SIZE-1) & MULT_95(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(19)(MULT_SIZE-1) & MULT_96(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(20)<=signed(MULT_95(20)(MULT_SIZE-1) & MULT_95(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(20)(MULT_SIZE-1) & MULT_96(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(21)<=signed(MULT_95(21)(MULT_SIZE-1) & MULT_95(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(21)(MULT_SIZE-1) & MULT_96(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(22)<=signed(MULT_95(22)(MULT_SIZE-1) & MULT_95(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(22)(MULT_SIZE-1) & MULT_96(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(23)<=signed(MULT_95(23)(MULT_SIZE-1) & MULT_95(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(23)(MULT_SIZE-1) & MULT_96(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(24)<=signed(MULT_95(24)(MULT_SIZE-1) & MULT_95(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(24)(MULT_SIZE-1) & MULT_96(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(25)<=signed(MULT_95(25)(MULT_SIZE-1) & MULT_95(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(25)(MULT_SIZE-1) & MULT_96(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(26)<=signed(MULT_95(26)(MULT_SIZE-1) & MULT_95(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(26)(MULT_SIZE-1) & MULT_96(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(27)<=signed(MULT_95(27)(MULT_SIZE-1) & MULT_95(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(27)(MULT_SIZE-1) & MULT_96(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(28)<=signed(MULT_95(28)(MULT_SIZE-1) & MULT_95(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(28)(MULT_SIZE-1) & MULT_96(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(29)<=signed(MULT_95(29)(MULT_SIZE-1) & MULT_95(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(29)(MULT_SIZE-1) & MULT_96(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(30)<=signed(MULT_95(30)(MULT_SIZE-1) & MULT_95(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(30)(MULT_SIZE-1) & MULT_96(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(31)<=signed(MULT_95(31)(MULT_SIZE-1) & MULT_95(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(31)(MULT_SIZE-1) & MULT_96(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(32)<=signed(MULT_95(32)(MULT_SIZE-1) & MULT_95(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(32)(MULT_SIZE-1) & MULT_96(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(33)<=signed(MULT_95(33)(MULT_SIZE-1) & MULT_95(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(33)(MULT_SIZE-1) & MULT_96(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(34)<=signed(MULT_95(34)(MULT_SIZE-1) & MULT_95(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(34)(MULT_SIZE-1) & MULT_96(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(35)<=signed(MULT_95(35)(MULT_SIZE-1) & MULT_95(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(35)(MULT_SIZE-1) & MULT_96(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(36)<=signed(MULT_95(36)(MULT_SIZE-1) & MULT_95(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(36)(MULT_SIZE-1) & MULT_96(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(37)<=signed(MULT_95(37)(MULT_SIZE-1) & MULT_95(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(37)(MULT_SIZE-1) & MULT_96(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(38)<=signed(MULT_95(38)(MULT_SIZE-1) & MULT_95(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(38)(MULT_SIZE-1) & MULT_96(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(39)<=signed(MULT_95(39)(MULT_SIZE-1) & MULT_95(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(39)(MULT_SIZE-1) & MULT_96(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(40)<=signed(MULT_95(40)(MULT_SIZE-1) & MULT_95(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(40)(MULT_SIZE-1) & MULT_96(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(41)<=signed(MULT_95(41)(MULT_SIZE-1) & MULT_95(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(41)(MULT_SIZE-1) & MULT_96(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(42)<=signed(MULT_95(42)(MULT_SIZE-1) & MULT_95(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(42)(MULT_SIZE-1) & MULT_96(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(43)<=signed(MULT_95(43)(MULT_SIZE-1) & MULT_95(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(43)(MULT_SIZE-1) & MULT_96(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(44)<=signed(MULT_95(44)(MULT_SIZE-1) & MULT_95(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(44)(MULT_SIZE-1) & MULT_96(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(45)<=signed(MULT_95(45)(MULT_SIZE-1) & MULT_95(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(45)(MULT_SIZE-1) & MULT_96(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(46)<=signed(MULT_95(46)(MULT_SIZE-1) & MULT_95(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(46)(MULT_SIZE-1) & MULT_96(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(47)<=signed(MULT_95(47)(MULT_SIZE-1) & MULT_95(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(47)(MULT_SIZE-1) & MULT_96(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(48)<=signed(MULT_95(48)(MULT_SIZE-1) & MULT_95(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(48)(MULT_SIZE-1) & MULT_96(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(49)<=signed(MULT_95(49)(MULT_SIZE-1) & MULT_95(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(49)(MULT_SIZE-1) & MULT_96(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(50)<=signed(MULT_95(50)(MULT_SIZE-1) & MULT_95(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(50)(MULT_SIZE-1) & MULT_96(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(51)<=signed(MULT_95(51)(MULT_SIZE-1) & MULT_95(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(51)(MULT_SIZE-1) & MULT_96(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(52)<=signed(MULT_95(52)(MULT_SIZE-1) & MULT_95(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(52)(MULT_SIZE-1) & MULT_96(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(53)<=signed(MULT_95(53)(MULT_SIZE-1) & MULT_95(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(53)(MULT_SIZE-1) & MULT_96(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(54)<=signed(MULT_95(54)(MULT_SIZE-1) & MULT_95(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(54)(MULT_SIZE-1) & MULT_96(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(55)<=signed(MULT_95(55)(MULT_SIZE-1) & MULT_95(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(55)(MULT_SIZE-1) & MULT_96(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(56)<=signed(MULT_95(56)(MULT_SIZE-1) & MULT_95(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(56)(MULT_SIZE-1) & MULT_96(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(57)<=signed(MULT_95(57)(MULT_SIZE-1) & MULT_95(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(57)(MULT_SIZE-1) & MULT_96(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(58)<=signed(MULT_95(58)(MULT_SIZE-1) & MULT_95(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(58)(MULT_SIZE-1) & MULT_96(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(59)<=signed(MULT_95(59)(MULT_SIZE-1) & MULT_95(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(59)(MULT_SIZE-1) & MULT_96(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(60)<=signed(MULT_95(60)(MULT_SIZE-1) & MULT_95(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(60)(MULT_SIZE-1) & MULT_96(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(61)<=signed(MULT_95(61)(MULT_SIZE-1) & MULT_95(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(61)(MULT_SIZE-1) & MULT_96(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(62)<=signed(MULT_95(62)(MULT_SIZE-1) & MULT_95(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(62)(MULT_SIZE-1) & MULT_96(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(63)<=signed(MULT_95(63)(MULT_SIZE-1) & MULT_95(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(63)(MULT_SIZE-1) & MULT_96(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(64)<=signed(MULT_95(64)(MULT_SIZE-1) & MULT_95(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(64)(MULT_SIZE-1) & MULT_96(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(65)<=signed(MULT_95(65)(MULT_SIZE-1) & MULT_95(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(65)(MULT_SIZE-1) & MULT_96(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(66)<=signed(MULT_95(66)(MULT_SIZE-1) & MULT_95(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(66)(MULT_SIZE-1) & MULT_96(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(67)<=signed(MULT_95(67)(MULT_SIZE-1) & MULT_95(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(67)(MULT_SIZE-1) & MULT_96(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(68)<=signed(MULT_95(68)(MULT_SIZE-1) & MULT_95(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(68)(MULT_SIZE-1) & MULT_96(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(69)<=signed(MULT_95(69)(MULT_SIZE-1) & MULT_95(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(69)(MULT_SIZE-1) & MULT_96(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(70)<=signed(MULT_95(70)(MULT_SIZE-1) & MULT_95(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(70)(MULT_SIZE-1) & MULT_96(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(71)<=signed(MULT_95(71)(MULT_SIZE-1) & MULT_95(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(71)(MULT_SIZE-1) & MULT_96(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(72)<=signed(MULT_95(72)(MULT_SIZE-1) & MULT_95(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(72)(MULT_SIZE-1) & MULT_96(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(73)<=signed(MULT_95(73)(MULT_SIZE-1) & MULT_95(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(73)(MULT_SIZE-1) & MULT_96(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(74)<=signed(MULT_95(74)(MULT_SIZE-1) & MULT_95(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(74)(MULT_SIZE-1) & MULT_96(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(75)<=signed(MULT_95(75)(MULT_SIZE-1) & MULT_95(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(75)(MULT_SIZE-1) & MULT_96(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(76)<=signed(MULT_95(76)(MULT_SIZE-1) & MULT_95(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(76)(MULT_SIZE-1) & MULT_96(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(77)<=signed(MULT_95(77)(MULT_SIZE-1) & MULT_95(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(77)(MULT_SIZE-1) & MULT_96(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(78)<=signed(MULT_95(78)(MULT_SIZE-1) & MULT_95(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(78)(MULT_SIZE-1) & MULT_96(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(79)<=signed(MULT_95(79)(MULT_SIZE-1) & MULT_95(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(79)(MULT_SIZE-1) & MULT_96(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(80)<=signed(MULT_95(80)(MULT_SIZE-1) & MULT_95(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(80)(MULT_SIZE-1) & MULT_96(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(81)<=signed(MULT_95(81)(MULT_SIZE-1) & MULT_95(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(81)(MULT_SIZE-1) & MULT_96(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(82)<=signed(MULT_95(82)(MULT_SIZE-1) & MULT_95(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(82)(MULT_SIZE-1) & MULT_96(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_48(83)<=signed(MULT_95(83)(MULT_SIZE-1) & MULT_95(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_96(83)(MULT_SIZE-1) & MULT_96(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_49(0)<=signed(MULT_97(0)(MULT_SIZE-1) & MULT_97(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(0)(MULT_SIZE-1) & MULT_98(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(1)<=signed(MULT_97(1)(MULT_SIZE-1) & MULT_97(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(1)(MULT_SIZE-1) & MULT_98(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(2)<=signed(MULT_97(2)(MULT_SIZE-1) & MULT_97(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(2)(MULT_SIZE-1) & MULT_98(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(3)<=signed(MULT_97(3)(MULT_SIZE-1) & MULT_97(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(3)(MULT_SIZE-1) & MULT_98(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(4)<=signed(MULT_97(4)(MULT_SIZE-1) & MULT_97(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(4)(MULT_SIZE-1) & MULT_98(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(5)<=signed(MULT_97(5)(MULT_SIZE-1) & MULT_97(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(5)(MULT_SIZE-1) & MULT_98(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(6)<=signed(MULT_97(6)(MULT_SIZE-1) & MULT_97(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(6)(MULT_SIZE-1) & MULT_98(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(7)<=signed(MULT_97(7)(MULT_SIZE-1) & MULT_97(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(7)(MULT_SIZE-1) & MULT_98(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(8)<=signed(MULT_97(8)(MULT_SIZE-1) & MULT_97(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(8)(MULT_SIZE-1) & MULT_98(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(9)<=signed(MULT_97(9)(MULT_SIZE-1) & MULT_97(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(9)(MULT_SIZE-1) & MULT_98(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(10)<=signed(MULT_97(10)(MULT_SIZE-1) & MULT_97(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(10)(MULT_SIZE-1) & MULT_98(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(11)<=signed(MULT_97(11)(MULT_SIZE-1) & MULT_97(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(11)(MULT_SIZE-1) & MULT_98(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(12)<=signed(MULT_97(12)(MULT_SIZE-1) & MULT_97(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(12)(MULT_SIZE-1) & MULT_98(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(13)<=signed(MULT_97(13)(MULT_SIZE-1) & MULT_97(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(13)(MULT_SIZE-1) & MULT_98(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(14)<=signed(MULT_97(14)(MULT_SIZE-1) & MULT_97(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(14)(MULT_SIZE-1) & MULT_98(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(15)<=signed(MULT_97(15)(MULT_SIZE-1) & MULT_97(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(15)(MULT_SIZE-1) & MULT_98(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(16)<=signed(MULT_97(16)(MULT_SIZE-1) & MULT_97(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(16)(MULT_SIZE-1) & MULT_98(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(17)<=signed(MULT_97(17)(MULT_SIZE-1) & MULT_97(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(17)(MULT_SIZE-1) & MULT_98(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(18)<=signed(MULT_97(18)(MULT_SIZE-1) & MULT_97(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(18)(MULT_SIZE-1) & MULT_98(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(19)<=signed(MULT_97(19)(MULT_SIZE-1) & MULT_97(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(19)(MULT_SIZE-1) & MULT_98(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(20)<=signed(MULT_97(20)(MULT_SIZE-1) & MULT_97(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(20)(MULT_SIZE-1) & MULT_98(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(21)<=signed(MULT_97(21)(MULT_SIZE-1) & MULT_97(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(21)(MULT_SIZE-1) & MULT_98(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(22)<=signed(MULT_97(22)(MULT_SIZE-1) & MULT_97(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(22)(MULT_SIZE-1) & MULT_98(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(23)<=signed(MULT_97(23)(MULT_SIZE-1) & MULT_97(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(23)(MULT_SIZE-1) & MULT_98(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(24)<=signed(MULT_97(24)(MULT_SIZE-1) & MULT_97(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(24)(MULT_SIZE-1) & MULT_98(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(25)<=signed(MULT_97(25)(MULT_SIZE-1) & MULT_97(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(25)(MULT_SIZE-1) & MULT_98(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(26)<=signed(MULT_97(26)(MULT_SIZE-1) & MULT_97(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(26)(MULT_SIZE-1) & MULT_98(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(27)<=signed(MULT_97(27)(MULT_SIZE-1) & MULT_97(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(27)(MULT_SIZE-1) & MULT_98(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(28)<=signed(MULT_97(28)(MULT_SIZE-1) & MULT_97(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(28)(MULT_SIZE-1) & MULT_98(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(29)<=signed(MULT_97(29)(MULT_SIZE-1) & MULT_97(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(29)(MULT_SIZE-1) & MULT_98(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(30)<=signed(MULT_97(30)(MULT_SIZE-1) & MULT_97(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(30)(MULT_SIZE-1) & MULT_98(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(31)<=signed(MULT_97(31)(MULT_SIZE-1) & MULT_97(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(31)(MULT_SIZE-1) & MULT_98(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(32)<=signed(MULT_97(32)(MULT_SIZE-1) & MULT_97(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(32)(MULT_SIZE-1) & MULT_98(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(33)<=signed(MULT_97(33)(MULT_SIZE-1) & MULT_97(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(33)(MULT_SIZE-1) & MULT_98(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(34)<=signed(MULT_97(34)(MULT_SIZE-1) & MULT_97(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(34)(MULT_SIZE-1) & MULT_98(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(35)<=signed(MULT_97(35)(MULT_SIZE-1) & MULT_97(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(35)(MULT_SIZE-1) & MULT_98(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(36)<=signed(MULT_97(36)(MULT_SIZE-1) & MULT_97(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(36)(MULT_SIZE-1) & MULT_98(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(37)<=signed(MULT_97(37)(MULT_SIZE-1) & MULT_97(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(37)(MULT_SIZE-1) & MULT_98(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(38)<=signed(MULT_97(38)(MULT_SIZE-1) & MULT_97(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(38)(MULT_SIZE-1) & MULT_98(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(39)<=signed(MULT_97(39)(MULT_SIZE-1) & MULT_97(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(39)(MULT_SIZE-1) & MULT_98(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(40)<=signed(MULT_97(40)(MULT_SIZE-1) & MULT_97(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(40)(MULT_SIZE-1) & MULT_98(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(41)<=signed(MULT_97(41)(MULT_SIZE-1) & MULT_97(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(41)(MULT_SIZE-1) & MULT_98(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(42)<=signed(MULT_97(42)(MULT_SIZE-1) & MULT_97(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(42)(MULT_SIZE-1) & MULT_98(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(43)<=signed(MULT_97(43)(MULT_SIZE-1) & MULT_97(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(43)(MULT_SIZE-1) & MULT_98(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(44)<=signed(MULT_97(44)(MULT_SIZE-1) & MULT_97(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(44)(MULT_SIZE-1) & MULT_98(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(45)<=signed(MULT_97(45)(MULT_SIZE-1) & MULT_97(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(45)(MULT_SIZE-1) & MULT_98(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(46)<=signed(MULT_97(46)(MULT_SIZE-1) & MULT_97(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(46)(MULT_SIZE-1) & MULT_98(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(47)<=signed(MULT_97(47)(MULT_SIZE-1) & MULT_97(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(47)(MULT_SIZE-1) & MULT_98(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(48)<=signed(MULT_97(48)(MULT_SIZE-1) & MULT_97(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(48)(MULT_SIZE-1) & MULT_98(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(49)<=signed(MULT_97(49)(MULT_SIZE-1) & MULT_97(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(49)(MULT_SIZE-1) & MULT_98(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(50)<=signed(MULT_97(50)(MULT_SIZE-1) & MULT_97(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(50)(MULT_SIZE-1) & MULT_98(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(51)<=signed(MULT_97(51)(MULT_SIZE-1) & MULT_97(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(51)(MULT_SIZE-1) & MULT_98(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(52)<=signed(MULT_97(52)(MULT_SIZE-1) & MULT_97(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(52)(MULT_SIZE-1) & MULT_98(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(53)<=signed(MULT_97(53)(MULT_SIZE-1) & MULT_97(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(53)(MULT_SIZE-1) & MULT_98(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(54)<=signed(MULT_97(54)(MULT_SIZE-1) & MULT_97(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(54)(MULT_SIZE-1) & MULT_98(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(55)<=signed(MULT_97(55)(MULT_SIZE-1) & MULT_97(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(55)(MULT_SIZE-1) & MULT_98(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(56)<=signed(MULT_97(56)(MULT_SIZE-1) & MULT_97(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(56)(MULT_SIZE-1) & MULT_98(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(57)<=signed(MULT_97(57)(MULT_SIZE-1) & MULT_97(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(57)(MULT_SIZE-1) & MULT_98(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(58)<=signed(MULT_97(58)(MULT_SIZE-1) & MULT_97(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(58)(MULT_SIZE-1) & MULT_98(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(59)<=signed(MULT_97(59)(MULT_SIZE-1) & MULT_97(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(59)(MULT_SIZE-1) & MULT_98(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(60)<=signed(MULT_97(60)(MULT_SIZE-1) & MULT_97(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(60)(MULT_SIZE-1) & MULT_98(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(61)<=signed(MULT_97(61)(MULT_SIZE-1) & MULT_97(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(61)(MULT_SIZE-1) & MULT_98(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(62)<=signed(MULT_97(62)(MULT_SIZE-1) & MULT_97(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(62)(MULT_SIZE-1) & MULT_98(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(63)<=signed(MULT_97(63)(MULT_SIZE-1) & MULT_97(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(63)(MULT_SIZE-1) & MULT_98(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(64)<=signed(MULT_97(64)(MULT_SIZE-1) & MULT_97(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(64)(MULT_SIZE-1) & MULT_98(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(65)<=signed(MULT_97(65)(MULT_SIZE-1) & MULT_97(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(65)(MULT_SIZE-1) & MULT_98(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(66)<=signed(MULT_97(66)(MULT_SIZE-1) & MULT_97(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(66)(MULT_SIZE-1) & MULT_98(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(67)<=signed(MULT_97(67)(MULT_SIZE-1) & MULT_97(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(67)(MULT_SIZE-1) & MULT_98(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(68)<=signed(MULT_97(68)(MULT_SIZE-1) & MULT_97(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(68)(MULT_SIZE-1) & MULT_98(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(69)<=signed(MULT_97(69)(MULT_SIZE-1) & MULT_97(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(69)(MULT_SIZE-1) & MULT_98(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(70)<=signed(MULT_97(70)(MULT_SIZE-1) & MULT_97(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(70)(MULT_SIZE-1) & MULT_98(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(71)<=signed(MULT_97(71)(MULT_SIZE-1) & MULT_97(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(71)(MULT_SIZE-1) & MULT_98(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(72)<=signed(MULT_97(72)(MULT_SIZE-1) & MULT_97(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(72)(MULT_SIZE-1) & MULT_98(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(73)<=signed(MULT_97(73)(MULT_SIZE-1) & MULT_97(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(73)(MULT_SIZE-1) & MULT_98(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(74)<=signed(MULT_97(74)(MULT_SIZE-1) & MULT_97(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(74)(MULT_SIZE-1) & MULT_98(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(75)<=signed(MULT_97(75)(MULT_SIZE-1) & MULT_97(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(75)(MULT_SIZE-1) & MULT_98(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(76)<=signed(MULT_97(76)(MULT_SIZE-1) & MULT_97(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(76)(MULT_SIZE-1) & MULT_98(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(77)<=signed(MULT_97(77)(MULT_SIZE-1) & MULT_97(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(77)(MULT_SIZE-1) & MULT_98(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(78)<=signed(MULT_97(78)(MULT_SIZE-1) & MULT_97(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(78)(MULT_SIZE-1) & MULT_98(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(79)<=signed(MULT_97(79)(MULT_SIZE-1) & MULT_97(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(79)(MULT_SIZE-1) & MULT_98(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(80)<=signed(MULT_97(80)(MULT_SIZE-1) & MULT_97(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(80)(MULT_SIZE-1) & MULT_98(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(81)<=signed(MULT_97(81)(MULT_SIZE-1) & MULT_97(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(81)(MULT_SIZE-1) & MULT_98(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(82)<=signed(MULT_97(82)(MULT_SIZE-1) & MULT_97(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(82)(MULT_SIZE-1) & MULT_98(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_49(83)<=signed(MULT_97(83)(MULT_SIZE-1) & MULT_97(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_98(83)(MULT_SIZE-1) & MULT_98(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_50(0)<=signed(MULT_99(0)(MULT_SIZE-1) & MULT_99(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(0)(MULT_SIZE-1) & MULT_100(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(1)<=signed(MULT_99(1)(MULT_SIZE-1) & MULT_99(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(1)(MULT_SIZE-1) & MULT_100(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(2)<=signed(MULT_99(2)(MULT_SIZE-1) & MULT_99(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(2)(MULT_SIZE-1) & MULT_100(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(3)<=signed(MULT_99(3)(MULT_SIZE-1) & MULT_99(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(3)(MULT_SIZE-1) & MULT_100(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(4)<=signed(MULT_99(4)(MULT_SIZE-1) & MULT_99(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(4)(MULT_SIZE-1) & MULT_100(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(5)<=signed(MULT_99(5)(MULT_SIZE-1) & MULT_99(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(5)(MULT_SIZE-1) & MULT_100(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(6)<=signed(MULT_99(6)(MULT_SIZE-1) & MULT_99(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(6)(MULT_SIZE-1) & MULT_100(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(7)<=signed(MULT_99(7)(MULT_SIZE-1) & MULT_99(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(7)(MULT_SIZE-1) & MULT_100(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(8)<=signed(MULT_99(8)(MULT_SIZE-1) & MULT_99(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(8)(MULT_SIZE-1) & MULT_100(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(9)<=signed(MULT_99(9)(MULT_SIZE-1) & MULT_99(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(9)(MULT_SIZE-1) & MULT_100(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(10)<=signed(MULT_99(10)(MULT_SIZE-1) & MULT_99(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(10)(MULT_SIZE-1) & MULT_100(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(11)<=signed(MULT_99(11)(MULT_SIZE-1) & MULT_99(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(11)(MULT_SIZE-1) & MULT_100(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(12)<=signed(MULT_99(12)(MULT_SIZE-1) & MULT_99(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(12)(MULT_SIZE-1) & MULT_100(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(13)<=signed(MULT_99(13)(MULT_SIZE-1) & MULT_99(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(13)(MULT_SIZE-1) & MULT_100(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(14)<=signed(MULT_99(14)(MULT_SIZE-1) & MULT_99(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(14)(MULT_SIZE-1) & MULT_100(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(15)<=signed(MULT_99(15)(MULT_SIZE-1) & MULT_99(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(15)(MULT_SIZE-1) & MULT_100(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(16)<=signed(MULT_99(16)(MULT_SIZE-1) & MULT_99(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(16)(MULT_SIZE-1) & MULT_100(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(17)<=signed(MULT_99(17)(MULT_SIZE-1) & MULT_99(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(17)(MULT_SIZE-1) & MULT_100(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(18)<=signed(MULT_99(18)(MULT_SIZE-1) & MULT_99(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(18)(MULT_SIZE-1) & MULT_100(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(19)<=signed(MULT_99(19)(MULT_SIZE-1) & MULT_99(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(19)(MULT_SIZE-1) & MULT_100(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(20)<=signed(MULT_99(20)(MULT_SIZE-1) & MULT_99(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(20)(MULT_SIZE-1) & MULT_100(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(21)<=signed(MULT_99(21)(MULT_SIZE-1) & MULT_99(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(21)(MULT_SIZE-1) & MULT_100(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(22)<=signed(MULT_99(22)(MULT_SIZE-1) & MULT_99(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(22)(MULT_SIZE-1) & MULT_100(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(23)<=signed(MULT_99(23)(MULT_SIZE-1) & MULT_99(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(23)(MULT_SIZE-1) & MULT_100(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(24)<=signed(MULT_99(24)(MULT_SIZE-1) & MULT_99(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(24)(MULT_SIZE-1) & MULT_100(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(25)<=signed(MULT_99(25)(MULT_SIZE-1) & MULT_99(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(25)(MULT_SIZE-1) & MULT_100(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(26)<=signed(MULT_99(26)(MULT_SIZE-1) & MULT_99(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(26)(MULT_SIZE-1) & MULT_100(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(27)<=signed(MULT_99(27)(MULT_SIZE-1) & MULT_99(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(27)(MULT_SIZE-1) & MULT_100(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(28)<=signed(MULT_99(28)(MULT_SIZE-1) & MULT_99(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(28)(MULT_SIZE-1) & MULT_100(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(29)<=signed(MULT_99(29)(MULT_SIZE-1) & MULT_99(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(29)(MULT_SIZE-1) & MULT_100(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(30)<=signed(MULT_99(30)(MULT_SIZE-1) & MULT_99(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(30)(MULT_SIZE-1) & MULT_100(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(31)<=signed(MULT_99(31)(MULT_SIZE-1) & MULT_99(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(31)(MULT_SIZE-1) & MULT_100(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(32)<=signed(MULT_99(32)(MULT_SIZE-1) & MULT_99(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(32)(MULT_SIZE-1) & MULT_100(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(33)<=signed(MULT_99(33)(MULT_SIZE-1) & MULT_99(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(33)(MULT_SIZE-1) & MULT_100(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(34)<=signed(MULT_99(34)(MULT_SIZE-1) & MULT_99(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(34)(MULT_SIZE-1) & MULT_100(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(35)<=signed(MULT_99(35)(MULT_SIZE-1) & MULT_99(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(35)(MULT_SIZE-1) & MULT_100(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(36)<=signed(MULT_99(36)(MULT_SIZE-1) & MULT_99(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(36)(MULT_SIZE-1) & MULT_100(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(37)<=signed(MULT_99(37)(MULT_SIZE-1) & MULT_99(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(37)(MULT_SIZE-1) & MULT_100(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(38)<=signed(MULT_99(38)(MULT_SIZE-1) & MULT_99(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(38)(MULT_SIZE-1) & MULT_100(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(39)<=signed(MULT_99(39)(MULT_SIZE-1) & MULT_99(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(39)(MULT_SIZE-1) & MULT_100(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(40)<=signed(MULT_99(40)(MULT_SIZE-1) & MULT_99(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(40)(MULT_SIZE-1) & MULT_100(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(41)<=signed(MULT_99(41)(MULT_SIZE-1) & MULT_99(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(41)(MULT_SIZE-1) & MULT_100(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(42)<=signed(MULT_99(42)(MULT_SIZE-1) & MULT_99(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(42)(MULT_SIZE-1) & MULT_100(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(43)<=signed(MULT_99(43)(MULT_SIZE-1) & MULT_99(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(43)(MULT_SIZE-1) & MULT_100(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(44)<=signed(MULT_99(44)(MULT_SIZE-1) & MULT_99(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(44)(MULT_SIZE-1) & MULT_100(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(45)<=signed(MULT_99(45)(MULT_SIZE-1) & MULT_99(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(45)(MULT_SIZE-1) & MULT_100(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(46)<=signed(MULT_99(46)(MULT_SIZE-1) & MULT_99(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(46)(MULT_SIZE-1) & MULT_100(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(47)<=signed(MULT_99(47)(MULT_SIZE-1) & MULT_99(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(47)(MULT_SIZE-1) & MULT_100(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(48)<=signed(MULT_99(48)(MULT_SIZE-1) & MULT_99(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(48)(MULT_SIZE-1) & MULT_100(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(49)<=signed(MULT_99(49)(MULT_SIZE-1) & MULT_99(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(49)(MULT_SIZE-1) & MULT_100(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(50)<=signed(MULT_99(50)(MULT_SIZE-1) & MULT_99(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(50)(MULT_SIZE-1) & MULT_100(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(51)<=signed(MULT_99(51)(MULT_SIZE-1) & MULT_99(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(51)(MULT_SIZE-1) & MULT_100(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(52)<=signed(MULT_99(52)(MULT_SIZE-1) & MULT_99(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(52)(MULT_SIZE-1) & MULT_100(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(53)<=signed(MULT_99(53)(MULT_SIZE-1) & MULT_99(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(53)(MULT_SIZE-1) & MULT_100(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(54)<=signed(MULT_99(54)(MULT_SIZE-1) & MULT_99(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(54)(MULT_SIZE-1) & MULT_100(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(55)<=signed(MULT_99(55)(MULT_SIZE-1) & MULT_99(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(55)(MULT_SIZE-1) & MULT_100(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(56)<=signed(MULT_99(56)(MULT_SIZE-1) & MULT_99(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(56)(MULT_SIZE-1) & MULT_100(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(57)<=signed(MULT_99(57)(MULT_SIZE-1) & MULT_99(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(57)(MULT_SIZE-1) & MULT_100(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(58)<=signed(MULT_99(58)(MULT_SIZE-1) & MULT_99(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(58)(MULT_SIZE-1) & MULT_100(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(59)<=signed(MULT_99(59)(MULT_SIZE-1) & MULT_99(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(59)(MULT_SIZE-1) & MULT_100(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(60)<=signed(MULT_99(60)(MULT_SIZE-1) & MULT_99(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(60)(MULT_SIZE-1) & MULT_100(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(61)<=signed(MULT_99(61)(MULT_SIZE-1) & MULT_99(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(61)(MULT_SIZE-1) & MULT_100(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(62)<=signed(MULT_99(62)(MULT_SIZE-1) & MULT_99(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(62)(MULT_SIZE-1) & MULT_100(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(63)<=signed(MULT_99(63)(MULT_SIZE-1) & MULT_99(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(63)(MULT_SIZE-1) & MULT_100(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(64)<=signed(MULT_99(64)(MULT_SIZE-1) & MULT_99(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(64)(MULT_SIZE-1) & MULT_100(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(65)<=signed(MULT_99(65)(MULT_SIZE-1) & MULT_99(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(65)(MULT_SIZE-1) & MULT_100(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(66)<=signed(MULT_99(66)(MULT_SIZE-1) & MULT_99(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(66)(MULT_SIZE-1) & MULT_100(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(67)<=signed(MULT_99(67)(MULT_SIZE-1) & MULT_99(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(67)(MULT_SIZE-1) & MULT_100(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(68)<=signed(MULT_99(68)(MULT_SIZE-1) & MULT_99(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(68)(MULT_SIZE-1) & MULT_100(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(69)<=signed(MULT_99(69)(MULT_SIZE-1) & MULT_99(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(69)(MULT_SIZE-1) & MULT_100(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(70)<=signed(MULT_99(70)(MULT_SIZE-1) & MULT_99(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(70)(MULT_SIZE-1) & MULT_100(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(71)<=signed(MULT_99(71)(MULT_SIZE-1) & MULT_99(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(71)(MULT_SIZE-1) & MULT_100(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(72)<=signed(MULT_99(72)(MULT_SIZE-1) & MULT_99(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(72)(MULT_SIZE-1) & MULT_100(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(73)<=signed(MULT_99(73)(MULT_SIZE-1) & MULT_99(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(73)(MULT_SIZE-1) & MULT_100(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(74)<=signed(MULT_99(74)(MULT_SIZE-1) & MULT_99(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(74)(MULT_SIZE-1) & MULT_100(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(75)<=signed(MULT_99(75)(MULT_SIZE-1) & MULT_99(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(75)(MULT_SIZE-1) & MULT_100(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(76)<=signed(MULT_99(76)(MULT_SIZE-1) & MULT_99(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(76)(MULT_SIZE-1) & MULT_100(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(77)<=signed(MULT_99(77)(MULT_SIZE-1) & MULT_99(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(77)(MULT_SIZE-1) & MULT_100(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(78)<=signed(MULT_99(78)(MULT_SIZE-1) & MULT_99(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(78)(MULT_SIZE-1) & MULT_100(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(79)<=signed(MULT_99(79)(MULT_SIZE-1) & MULT_99(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(79)(MULT_SIZE-1) & MULT_100(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(80)<=signed(MULT_99(80)(MULT_SIZE-1) & MULT_99(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(80)(MULT_SIZE-1) & MULT_100(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(81)<=signed(MULT_99(81)(MULT_SIZE-1) & MULT_99(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(81)(MULT_SIZE-1) & MULT_100(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(82)<=signed(MULT_99(82)(MULT_SIZE-1) & MULT_99(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(82)(MULT_SIZE-1) & MULT_100(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_50(83)<=signed(MULT_99(83)(MULT_SIZE-1) & MULT_99(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_100(83)(MULT_SIZE-1) & MULT_100(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_51(0)<=signed(MULT_101(0)(MULT_SIZE-1) & MULT_101(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(0)(MULT_SIZE-1) & MULT_102(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(1)<=signed(MULT_101(1)(MULT_SIZE-1) & MULT_101(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(1)(MULT_SIZE-1) & MULT_102(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(2)<=signed(MULT_101(2)(MULT_SIZE-1) & MULT_101(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(2)(MULT_SIZE-1) & MULT_102(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(3)<=signed(MULT_101(3)(MULT_SIZE-1) & MULT_101(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(3)(MULT_SIZE-1) & MULT_102(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(4)<=signed(MULT_101(4)(MULT_SIZE-1) & MULT_101(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(4)(MULT_SIZE-1) & MULT_102(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(5)<=signed(MULT_101(5)(MULT_SIZE-1) & MULT_101(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(5)(MULT_SIZE-1) & MULT_102(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(6)<=signed(MULT_101(6)(MULT_SIZE-1) & MULT_101(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(6)(MULT_SIZE-1) & MULT_102(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(7)<=signed(MULT_101(7)(MULT_SIZE-1) & MULT_101(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(7)(MULT_SIZE-1) & MULT_102(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(8)<=signed(MULT_101(8)(MULT_SIZE-1) & MULT_101(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(8)(MULT_SIZE-1) & MULT_102(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(9)<=signed(MULT_101(9)(MULT_SIZE-1) & MULT_101(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(9)(MULT_SIZE-1) & MULT_102(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(10)<=signed(MULT_101(10)(MULT_SIZE-1) & MULT_101(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(10)(MULT_SIZE-1) & MULT_102(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(11)<=signed(MULT_101(11)(MULT_SIZE-1) & MULT_101(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(11)(MULT_SIZE-1) & MULT_102(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(12)<=signed(MULT_101(12)(MULT_SIZE-1) & MULT_101(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(12)(MULT_SIZE-1) & MULT_102(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(13)<=signed(MULT_101(13)(MULT_SIZE-1) & MULT_101(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(13)(MULT_SIZE-1) & MULT_102(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(14)<=signed(MULT_101(14)(MULT_SIZE-1) & MULT_101(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(14)(MULT_SIZE-1) & MULT_102(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(15)<=signed(MULT_101(15)(MULT_SIZE-1) & MULT_101(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(15)(MULT_SIZE-1) & MULT_102(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(16)<=signed(MULT_101(16)(MULT_SIZE-1) & MULT_101(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(16)(MULT_SIZE-1) & MULT_102(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(17)<=signed(MULT_101(17)(MULT_SIZE-1) & MULT_101(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(17)(MULT_SIZE-1) & MULT_102(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(18)<=signed(MULT_101(18)(MULT_SIZE-1) & MULT_101(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(18)(MULT_SIZE-1) & MULT_102(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(19)<=signed(MULT_101(19)(MULT_SIZE-1) & MULT_101(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(19)(MULT_SIZE-1) & MULT_102(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(20)<=signed(MULT_101(20)(MULT_SIZE-1) & MULT_101(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(20)(MULT_SIZE-1) & MULT_102(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(21)<=signed(MULT_101(21)(MULT_SIZE-1) & MULT_101(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(21)(MULT_SIZE-1) & MULT_102(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(22)<=signed(MULT_101(22)(MULT_SIZE-1) & MULT_101(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(22)(MULT_SIZE-1) & MULT_102(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(23)<=signed(MULT_101(23)(MULT_SIZE-1) & MULT_101(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(23)(MULT_SIZE-1) & MULT_102(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(24)<=signed(MULT_101(24)(MULT_SIZE-1) & MULT_101(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(24)(MULT_SIZE-1) & MULT_102(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(25)<=signed(MULT_101(25)(MULT_SIZE-1) & MULT_101(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(25)(MULT_SIZE-1) & MULT_102(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(26)<=signed(MULT_101(26)(MULT_SIZE-1) & MULT_101(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(26)(MULT_SIZE-1) & MULT_102(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(27)<=signed(MULT_101(27)(MULT_SIZE-1) & MULT_101(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(27)(MULT_SIZE-1) & MULT_102(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(28)<=signed(MULT_101(28)(MULT_SIZE-1) & MULT_101(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(28)(MULT_SIZE-1) & MULT_102(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(29)<=signed(MULT_101(29)(MULT_SIZE-1) & MULT_101(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(29)(MULT_SIZE-1) & MULT_102(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(30)<=signed(MULT_101(30)(MULT_SIZE-1) & MULT_101(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(30)(MULT_SIZE-1) & MULT_102(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(31)<=signed(MULT_101(31)(MULT_SIZE-1) & MULT_101(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(31)(MULT_SIZE-1) & MULT_102(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(32)<=signed(MULT_101(32)(MULT_SIZE-1) & MULT_101(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(32)(MULT_SIZE-1) & MULT_102(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(33)<=signed(MULT_101(33)(MULT_SIZE-1) & MULT_101(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(33)(MULT_SIZE-1) & MULT_102(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(34)<=signed(MULT_101(34)(MULT_SIZE-1) & MULT_101(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(34)(MULT_SIZE-1) & MULT_102(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(35)<=signed(MULT_101(35)(MULT_SIZE-1) & MULT_101(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(35)(MULT_SIZE-1) & MULT_102(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(36)<=signed(MULT_101(36)(MULT_SIZE-1) & MULT_101(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(36)(MULT_SIZE-1) & MULT_102(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(37)<=signed(MULT_101(37)(MULT_SIZE-1) & MULT_101(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(37)(MULT_SIZE-1) & MULT_102(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(38)<=signed(MULT_101(38)(MULT_SIZE-1) & MULT_101(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(38)(MULT_SIZE-1) & MULT_102(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(39)<=signed(MULT_101(39)(MULT_SIZE-1) & MULT_101(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(39)(MULT_SIZE-1) & MULT_102(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(40)<=signed(MULT_101(40)(MULT_SIZE-1) & MULT_101(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(40)(MULT_SIZE-1) & MULT_102(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(41)<=signed(MULT_101(41)(MULT_SIZE-1) & MULT_101(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(41)(MULT_SIZE-1) & MULT_102(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(42)<=signed(MULT_101(42)(MULT_SIZE-1) & MULT_101(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(42)(MULT_SIZE-1) & MULT_102(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(43)<=signed(MULT_101(43)(MULT_SIZE-1) & MULT_101(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(43)(MULT_SIZE-1) & MULT_102(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(44)<=signed(MULT_101(44)(MULT_SIZE-1) & MULT_101(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(44)(MULT_SIZE-1) & MULT_102(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(45)<=signed(MULT_101(45)(MULT_SIZE-1) & MULT_101(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(45)(MULT_SIZE-1) & MULT_102(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(46)<=signed(MULT_101(46)(MULT_SIZE-1) & MULT_101(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(46)(MULT_SIZE-1) & MULT_102(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(47)<=signed(MULT_101(47)(MULT_SIZE-1) & MULT_101(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(47)(MULT_SIZE-1) & MULT_102(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(48)<=signed(MULT_101(48)(MULT_SIZE-1) & MULT_101(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(48)(MULT_SIZE-1) & MULT_102(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(49)<=signed(MULT_101(49)(MULT_SIZE-1) & MULT_101(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(49)(MULT_SIZE-1) & MULT_102(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(50)<=signed(MULT_101(50)(MULT_SIZE-1) & MULT_101(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(50)(MULT_SIZE-1) & MULT_102(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(51)<=signed(MULT_101(51)(MULT_SIZE-1) & MULT_101(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(51)(MULT_SIZE-1) & MULT_102(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(52)<=signed(MULT_101(52)(MULT_SIZE-1) & MULT_101(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(52)(MULT_SIZE-1) & MULT_102(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(53)<=signed(MULT_101(53)(MULT_SIZE-1) & MULT_101(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(53)(MULT_SIZE-1) & MULT_102(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(54)<=signed(MULT_101(54)(MULT_SIZE-1) & MULT_101(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(54)(MULT_SIZE-1) & MULT_102(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(55)<=signed(MULT_101(55)(MULT_SIZE-1) & MULT_101(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(55)(MULT_SIZE-1) & MULT_102(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(56)<=signed(MULT_101(56)(MULT_SIZE-1) & MULT_101(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(56)(MULT_SIZE-1) & MULT_102(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(57)<=signed(MULT_101(57)(MULT_SIZE-1) & MULT_101(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(57)(MULT_SIZE-1) & MULT_102(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(58)<=signed(MULT_101(58)(MULT_SIZE-1) & MULT_101(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(58)(MULT_SIZE-1) & MULT_102(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(59)<=signed(MULT_101(59)(MULT_SIZE-1) & MULT_101(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(59)(MULT_SIZE-1) & MULT_102(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(60)<=signed(MULT_101(60)(MULT_SIZE-1) & MULT_101(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(60)(MULT_SIZE-1) & MULT_102(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(61)<=signed(MULT_101(61)(MULT_SIZE-1) & MULT_101(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(61)(MULT_SIZE-1) & MULT_102(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(62)<=signed(MULT_101(62)(MULT_SIZE-1) & MULT_101(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(62)(MULT_SIZE-1) & MULT_102(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(63)<=signed(MULT_101(63)(MULT_SIZE-1) & MULT_101(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(63)(MULT_SIZE-1) & MULT_102(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(64)<=signed(MULT_101(64)(MULT_SIZE-1) & MULT_101(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(64)(MULT_SIZE-1) & MULT_102(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(65)<=signed(MULT_101(65)(MULT_SIZE-1) & MULT_101(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(65)(MULT_SIZE-1) & MULT_102(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(66)<=signed(MULT_101(66)(MULT_SIZE-1) & MULT_101(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(66)(MULT_SIZE-1) & MULT_102(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(67)<=signed(MULT_101(67)(MULT_SIZE-1) & MULT_101(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(67)(MULT_SIZE-1) & MULT_102(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(68)<=signed(MULT_101(68)(MULT_SIZE-1) & MULT_101(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(68)(MULT_SIZE-1) & MULT_102(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(69)<=signed(MULT_101(69)(MULT_SIZE-1) & MULT_101(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(69)(MULT_SIZE-1) & MULT_102(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(70)<=signed(MULT_101(70)(MULT_SIZE-1) & MULT_101(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(70)(MULT_SIZE-1) & MULT_102(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(71)<=signed(MULT_101(71)(MULT_SIZE-1) & MULT_101(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(71)(MULT_SIZE-1) & MULT_102(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(72)<=signed(MULT_101(72)(MULT_SIZE-1) & MULT_101(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(72)(MULT_SIZE-1) & MULT_102(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(73)<=signed(MULT_101(73)(MULT_SIZE-1) & MULT_101(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(73)(MULT_SIZE-1) & MULT_102(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(74)<=signed(MULT_101(74)(MULT_SIZE-1) & MULT_101(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(74)(MULT_SIZE-1) & MULT_102(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(75)<=signed(MULT_101(75)(MULT_SIZE-1) & MULT_101(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(75)(MULT_SIZE-1) & MULT_102(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(76)<=signed(MULT_101(76)(MULT_SIZE-1) & MULT_101(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(76)(MULT_SIZE-1) & MULT_102(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(77)<=signed(MULT_101(77)(MULT_SIZE-1) & MULT_101(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(77)(MULT_SIZE-1) & MULT_102(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(78)<=signed(MULT_101(78)(MULT_SIZE-1) & MULT_101(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(78)(MULT_SIZE-1) & MULT_102(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(79)<=signed(MULT_101(79)(MULT_SIZE-1) & MULT_101(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(79)(MULT_SIZE-1) & MULT_102(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(80)<=signed(MULT_101(80)(MULT_SIZE-1) & MULT_101(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(80)(MULT_SIZE-1) & MULT_102(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(81)<=signed(MULT_101(81)(MULT_SIZE-1) & MULT_101(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(81)(MULT_SIZE-1) & MULT_102(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(82)<=signed(MULT_101(82)(MULT_SIZE-1) & MULT_101(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(82)(MULT_SIZE-1) & MULT_102(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_51(83)<=signed(MULT_101(83)(MULT_SIZE-1) & MULT_101(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_102(83)(MULT_SIZE-1) & MULT_102(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_52(0)<=signed(MULT_103(0)(MULT_SIZE-1) & MULT_103(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(0)(MULT_SIZE-1) & MULT_104(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(1)<=signed(MULT_103(1)(MULT_SIZE-1) & MULT_103(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(1)(MULT_SIZE-1) & MULT_104(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(2)<=signed(MULT_103(2)(MULT_SIZE-1) & MULT_103(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(2)(MULT_SIZE-1) & MULT_104(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(3)<=signed(MULT_103(3)(MULT_SIZE-1) & MULT_103(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(3)(MULT_SIZE-1) & MULT_104(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(4)<=signed(MULT_103(4)(MULT_SIZE-1) & MULT_103(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(4)(MULT_SIZE-1) & MULT_104(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(5)<=signed(MULT_103(5)(MULT_SIZE-1) & MULT_103(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(5)(MULT_SIZE-1) & MULT_104(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(6)<=signed(MULT_103(6)(MULT_SIZE-1) & MULT_103(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(6)(MULT_SIZE-1) & MULT_104(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(7)<=signed(MULT_103(7)(MULT_SIZE-1) & MULT_103(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(7)(MULT_SIZE-1) & MULT_104(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(8)<=signed(MULT_103(8)(MULT_SIZE-1) & MULT_103(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(8)(MULT_SIZE-1) & MULT_104(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(9)<=signed(MULT_103(9)(MULT_SIZE-1) & MULT_103(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(9)(MULT_SIZE-1) & MULT_104(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(10)<=signed(MULT_103(10)(MULT_SIZE-1) & MULT_103(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(10)(MULT_SIZE-1) & MULT_104(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(11)<=signed(MULT_103(11)(MULT_SIZE-1) & MULT_103(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(11)(MULT_SIZE-1) & MULT_104(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(12)<=signed(MULT_103(12)(MULT_SIZE-1) & MULT_103(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(12)(MULT_SIZE-1) & MULT_104(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(13)<=signed(MULT_103(13)(MULT_SIZE-1) & MULT_103(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(13)(MULT_SIZE-1) & MULT_104(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(14)<=signed(MULT_103(14)(MULT_SIZE-1) & MULT_103(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(14)(MULT_SIZE-1) & MULT_104(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(15)<=signed(MULT_103(15)(MULT_SIZE-1) & MULT_103(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(15)(MULT_SIZE-1) & MULT_104(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(16)<=signed(MULT_103(16)(MULT_SIZE-1) & MULT_103(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(16)(MULT_SIZE-1) & MULT_104(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(17)<=signed(MULT_103(17)(MULT_SIZE-1) & MULT_103(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(17)(MULT_SIZE-1) & MULT_104(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(18)<=signed(MULT_103(18)(MULT_SIZE-1) & MULT_103(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(18)(MULT_SIZE-1) & MULT_104(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(19)<=signed(MULT_103(19)(MULT_SIZE-1) & MULT_103(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(19)(MULT_SIZE-1) & MULT_104(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(20)<=signed(MULT_103(20)(MULT_SIZE-1) & MULT_103(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(20)(MULT_SIZE-1) & MULT_104(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(21)<=signed(MULT_103(21)(MULT_SIZE-1) & MULT_103(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(21)(MULT_SIZE-1) & MULT_104(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(22)<=signed(MULT_103(22)(MULT_SIZE-1) & MULT_103(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(22)(MULT_SIZE-1) & MULT_104(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(23)<=signed(MULT_103(23)(MULT_SIZE-1) & MULT_103(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(23)(MULT_SIZE-1) & MULT_104(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(24)<=signed(MULT_103(24)(MULT_SIZE-1) & MULT_103(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(24)(MULT_SIZE-1) & MULT_104(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(25)<=signed(MULT_103(25)(MULT_SIZE-1) & MULT_103(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(25)(MULT_SIZE-1) & MULT_104(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(26)<=signed(MULT_103(26)(MULT_SIZE-1) & MULT_103(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(26)(MULT_SIZE-1) & MULT_104(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(27)<=signed(MULT_103(27)(MULT_SIZE-1) & MULT_103(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(27)(MULT_SIZE-1) & MULT_104(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(28)<=signed(MULT_103(28)(MULT_SIZE-1) & MULT_103(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(28)(MULT_SIZE-1) & MULT_104(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(29)<=signed(MULT_103(29)(MULT_SIZE-1) & MULT_103(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(29)(MULT_SIZE-1) & MULT_104(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(30)<=signed(MULT_103(30)(MULT_SIZE-1) & MULT_103(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(30)(MULT_SIZE-1) & MULT_104(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(31)<=signed(MULT_103(31)(MULT_SIZE-1) & MULT_103(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(31)(MULT_SIZE-1) & MULT_104(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(32)<=signed(MULT_103(32)(MULT_SIZE-1) & MULT_103(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(32)(MULT_SIZE-1) & MULT_104(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(33)<=signed(MULT_103(33)(MULT_SIZE-1) & MULT_103(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(33)(MULT_SIZE-1) & MULT_104(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(34)<=signed(MULT_103(34)(MULT_SIZE-1) & MULT_103(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(34)(MULT_SIZE-1) & MULT_104(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(35)<=signed(MULT_103(35)(MULT_SIZE-1) & MULT_103(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(35)(MULT_SIZE-1) & MULT_104(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(36)<=signed(MULT_103(36)(MULT_SIZE-1) & MULT_103(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(36)(MULT_SIZE-1) & MULT_104(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(37)<=signed(MULT_103(37)(MULT_SIZE-1) & MULT_103(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(37)(MULT_SIZE-1) & MULT_104(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(38)<=signed(MULT_103(38)(MULT_SIZE-1) & MULT_103(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(38)(MULT_SIZE-1) & MULT_104(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(39)<=signed(MULT_103(39)(MULT_SIZE-1) & MULT_103(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(39)(MULT_SIZE-1) & MULT_104(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(40)<=signed(MULT_103(40)(MULT_SIZE-1) & MULT_103(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(40)(MULT_SIZE-1) & MULT_104(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(41)<=signed(MULT_103(41)(MULT_SIZE-1) & MULT_103(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(41)(MULT_SIZE-1) & MULT_104(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(42)<=signed(MULT_103(42)(MULT_SIZE-1) & MULT_103(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(42)(MULT_SIZE-1) & MULT_104(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(43)<=signed(MULT_103(43)(MULT_SIZE-1) & MULT_103(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(43)(MULT_SIZE-1) & MULT_104(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(44)<=signed(MULT_103(44)(MULT_SIZE-1) & MULT_103(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(44)(MULT_SIZE-1) & MULT_104(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(45)<=signed(MULT_103(45)(MULT_SIZE-1) & MULT_103(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(45)(MULT_SIZE-1) & MULT_104(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(46)<=signed(MULT_103(46)(MULT_SIZE-1) & MULT_103(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(46)(MULT_SIZE-1) & MULT_104(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(47)<=signed(MULT_103(47)(MULT_SIZE-1) & MULT_103(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(47)(MULT_SIZE-1) & MULT_104(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(48)<=signed(MULT_103(48)(MULT_SIZE-1) & MULT_103(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(48)(MULT_SIZE-1) & MULT_104(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(49)<=signed(MULT_103(49)(MULT_SIZE-1) & MULT_103(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(49)(MULT_SIZE-1) & MULT_104(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(50)<=signed(MULT_103(50)(MULT_SIZE-1) & MULT_103(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(50)(MULT_SIZE-1) & MULT_104(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(51)<=signed(MULT_103(51)(MULT_SIZE-1) & MULT_103(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(51)(MULT_SIZE-1) & MULT_104(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(52)<=signed(MULT_103(52)(MULT_SIZE-1) & MULT_103(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(52)(MULT_SIZE-1) & MULT_104(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(53)<=signed(MULT_103(53)(MULT_SIZE-1) & MULT_103(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(53)(MULT_SIZE-1) & MULT_104(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(54)<=signed(MULT_103(54)(MULT_SIZE-1) & MULT_103(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(54)(MULT_SIZE-1) & MULT_104(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(55)<=signed(MULT_103(55)(MULT_SIZE-1) & MULT_103(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(55)(MULT_SIZE-1) & MULT_104(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(56)<=signed(MULT_103(56)(MULT_SIZE-1) & MULT_103(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(56)(MULT_SIZE-1) & MULT_104(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(57)<=signed(MULT_103(57)(MULT_SIZE-1) & MULT_103(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(57)(MULT_SIZE-1) & MULT_104(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(58)<=signed(MULT_103(58)(MULT_SIZE-1) & MULT_103(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(58)(MULT_SIZE-1) & MULT_104(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(59)<=signed(MULT_103(59)(MULT_SIZE-1) & MULT_103(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(59)(MULT_SIZE-1) & MULT_104(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(60)<=signed(MULT_103(60)(MULT_SIZE-1) & MULT_103(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(60)(MULT_SIZE-1) & MULT_104(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(61)<=signed(MULT_103(61)(MULT_SIZE-1) & MULT_103(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(61)(MULT_SIZE-1) & MULT_104(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(62)<=signed(MULT_103(62)(MULT_SIZE-1) & MULT_103(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(62)(MULT_SIZE-1) & MULT_104(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(63)<=signed(MULT_103(63)(MULT_SIZE-1) & MULT_103(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(63)(MULT_SIZE-1) & MULT_104(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(64)<=signed(MULT_103(64)(MULT_SIZE-1) & MULT_103(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(64)(MULT_SIZE-1) & MULT_104(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(65)<=signed(MULT_103(65)(MULT_SIZE-1) & MULT_103(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(65)(MULT_SIZE-1) & MULT_104(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(66)<=signed(MULT_103(66)(MULT_SIZE-1) & MULT_103(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(66)(MULT_SIZE-1) & MULT_104(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(67)<=signed(MULT_103(67)(MULT_SIZE-1) & MULT_103(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(67)(MULT_SIZE-1) & MULT_104(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(68)<=signed(MULT_103(68)(MULT_SIZE-1) & MULT_103(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(68)(MULT_SIZE-1) & MULT_104(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(69)<=signed(MULT_103(69)(MULT_SIZE-1) & MULT_103(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(69)(MULT_SIZE-1) & MULT_104(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(70)<=signed(MULT_103(70)(MULT_SIZE-1) & MULT_103(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(70)(MULT_SIZE-1) & MULT_104(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(71)<=signed(MULT_103(71)(MULT_SIZE-1) & MULT_103(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(71)(MULT_SIZE-1) & MULT_104(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(72)<=signed(MULT_103(72)(MULT_SIZE-1) & MULT_103(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(72)(MULT_SIZE-1) & MULT_104(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(73)<=signed(MULT_103(73)(MULT_SIZE-1) & MULT_103(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(73)(MULT_SIZE-1) & MULT_104(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(74)<=signed(MULT_103(74)(MULT_SIZE-1) & MULT_103(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(74)(MULT_SIZE-1) & MULT_104(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(75)<=signed(MULT_103(75)(MULT_SIZE-1) & MULT_103(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(75)(MULT_SIZE-1) & MULT_104(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(76)<=signed(MULT_103(76)(MULT_SIZE-1) & MULT_103(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(76)(MULT_SIZE-1) & MULT_104(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(77)<=signed(MULT_103(77)(MULT_SIZE-1) & MULT_103(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(77)(MULT_SIZE-1) & MULT_104(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(78)<=signed(MULT_103(78)(MULT_SIZE-1) & MULT_103(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(78)(MULT_SIZE-1) & MULT_104(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(79)<=signed(MULT_103(79)(MULT_SIZE-1) & MULT_103(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(79)(MULT_SIZE-1) & MULT_104(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(80)<=signed(MULT_103(80)(MULT_SIZE-1) & MULT_103(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(80)(MULT_SIZE-1) & MULT_104(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(81)<=signed(MULT_103(81)(MULT_SIZE-1) & MULT_103(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(81)(MULT_SIZE-1) & MULT_104(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(82)<=signed(MULT_103(82)(MULT_SIZE-1) & MULT_103(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(82)(MULT_SIZE-1) & MULT_104(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_52(83)<=signed(MULT_103(83)(MULT_SIZE-1) & MULT_103(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_104(83)(MULT_SIZE-1) & MULT_104(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_53(0)<=signed(MULT_105(0)(MULT_SIZE-1) & MULT_105(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(0)(MULT_SIZE-1) & MULT_106(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(1)<=signed(MULT_105(1)(MULT_SIZE-1) & MULT_105(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(1)(MULT_SIZE-1) & MULT_106(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(2)<=signed(MULT_105(2)(MULT_SIZE-1) & MULT_105(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(2)(MULT_SIZE-1) & MULT_106(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(3)<=signed(MULT_105(3)(MULT_SIZE-1) & MULT_105(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(3)(MULT_SIZE-1) & MULT_106(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(4)<=signed(MULT_105(4)(MULT_SIZE-1) & MULT_105(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(4)(MULT_SIZE-1) & MULT_106(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(5)<=signed(MULT_105(5)(MULT_SIZE-1) & MULT_105(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(5)(MULT_SIZE-1) & MULT_106(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(6)<=signed(MULT_105(6)(MULT_SIZE-1) & MULT_105(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(6)(MULT_SIZE-1) & MULT_106(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(7)<=signed(MULT_105(7)(MULT_SIZE-1) & MULT_105(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(7)(MULT_SIZE-1) & MULT_106(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(8)<=signed(MULT_105(8)(MULT_SIZE-1) & MULT_105(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(8)(MULT_SIZE-1) & MULT_106(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(9)<=signed(MULT_105(9)(MULT_SIZE-1) & MULT_105(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(9)(MULT_SIZE-1) & MULT_106(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(10)<=signed(MULT_105(10)(MULT_SIZE-1) & MULT_105(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(10)(MULT_SIZE-1) & MULT_106(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(11)<=signed(MULT_105(11)(MULT_SIZE-1) & MULT_105(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(11)(MULT_SIZE-1) & MULT_106(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(12)<=signed(MULT_105(12)(MULT_SIZE-1) & MULT_105(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(12)(MULT_SIZE-1) & MULT_106(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(13)<=signed(MULT_105(13)(MULT_SIZE-1) & MULT_105(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(13)(MULT_SIZE-1) & MULT_106(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(14)<=signed(MULT_105(14)(MULT_SIZE-1) & MULT_105(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(14)(MULT_SIZE-1) & MULT_106(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(15)<=signed(MULT_105(15)(MULT_SIZE-1) & MULT_105(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(15)(MULT_SIZE-1) & MULT_106(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(16)<=signed(MULT_105(16)(MULT_SIZE-1) & MULT_105(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(16)(MULT_SIZE-1) & MULT_106(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(17)<=signed(MULT_105(17)(MULT_SIZE-1) & MULT_105(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(17)(MULT_SIZE-1) & MULT_106(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(18)<=signed(MULT_105(18)(MULT_SIZE-1) & MULT_105(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(18)(MULT_SIZE-1) & MULT_106(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(19)<=signed(MULT_105(19)(MULT_SIZE-1) & MULT_105(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(19)(MULT_SIZE-1) & MULT_106(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(20)<=signed(MULT_105(20)(MULT_SIZE-1) & MULT_105(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(20)(MULT_SIZE-1) & MULT_106(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(21)<=signed(MULT_105(21)(MULT_SIZE-1) & MULT_105(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(21)(MULT_SIZE-1) & MULT_106(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(22)<=signed(MULT_105(22)(MULT_SIZE-1) & MULT_105(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(22)(MULT_SIZE-1) & MULT_106(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(23)<=signed(MULT_105(23)(MULT_SIZE-1) & MULT_105(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(23)(MULT_SIZE-1) & MULT_106(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(24)<=signed(MULT_105(24)(MULT_SIZE-1) & MULT_105(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(24)(MULT_SIZE-1) & MULT_106(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(25)<=signed(MULT_105(25)(MULT_SIZE-1) & MULT_105(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(25)(MULT_SIZE-1) & MULT_106(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(26)<=signed(MULT_105(26)(MULT_SIZE-1) & MULT_105(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(26)(MULT_SIZE-1) & MULT_106(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(27)<=signed(MULT_105(27)(MULT_SIZE-1) & MULT_105(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(27)(MULT_SIZE-1) & MULT_106(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(28)<=signed(MULT_105(28)(MULT_SIZE-1) & MULT_105(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(28)(MULT_SIZE-1) & MULT_106(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(29)<=signed(MULT_105(29)(MULT_SIZE-1) & MULT_105(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(29)(MULT_SIZE-1) & MULT_106(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(30)<=signed(MULT_105(30)(MULT_SIZE-1) & MULT_105(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(30)(MULT_SIZE-1) & MULT_106(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(31)<=signed(MULT_105(31)(MULT_SIZE-1) & MULT_105(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(31)(MULT_SIZE-1) & MULT_106(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(32)<=signed(MULT_105(32)(MULT_SIZE-1) & MULT_105(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(32)(MULT_SIZE-1) & MULT_106(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(33)<=signed(MULT_105(33)(MULT_SIZE-1) & MULT_105(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(33)(MULT_SIZE-1) & MULT_106(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(34)<=signed(MULT_105(34)(MULT_SIZE-1) & MULT_105(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(34)(MULT_SIZE-1) & MULT_106(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(35)<=signed(MULT_105(35)(MULT_SIZE-1) & MULT_105(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(35)(MULT_SIZE-1) & MULT_106(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(36)<=signed(MULT_105(36)(MULT_SIZE-1) & MULT_105(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(36)(MULT_SIZE-1) & MULT_106(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(37)<=signed(MULT_105(37)(MULT_SIZE-1) & MULT_105(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(37)(MULT_SIZE-1) & MULT_106(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(38)<=signed(MULT_105(38)(MULT_SIZE-1) & MULT_105(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(38)(MULT_SIZE-1) & MULT_106(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(39)<=signed(MULT_105(39)(MULT_SIZE-1) & MULT_105(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(39)(MULT_SIZE-1) & MULT_106(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(40)<=signed(MULT_105(40)(MULT_SIZE-1) & MULT_105(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(40)(MULT_SIZE-1) & MULT_106(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(41)<=signed(MULT_105(41)(MULT_SIZE-1) & MULT_105(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(41)(MULT_SIZE-1) & MULT_106(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(42)<=signed(MULT_105(42)(MULT_SIZE-1) & MULT_105(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(42)(MULT_SIZE-1) & MULT_106(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(43)<=signed(MULT_105(43)(MULT_SIZE-1) & MULT_105(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(43)(MULT_SIZE-1) & MULT_106(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(44)<=signed(MULT_105(44)(MULT_SIZE-1) & MULT_105(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(44)(MULT_SIZE-1) & MULT_106(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(45)<=signed(MULT_105(45)(MULT_SIZE-1) & MULT_105(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(45)(MULT_SIZE-1) & MULT_106(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(46)<=signed(MULT_105(46)(MULT_SIZE-1) & MULT_105(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(46)(MULT_SIZE-1) & MULT_106(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(47)<=signed(MULT_105(47)(MULT_SIZE-1) & MULT_105(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(47)(MULT_SIZE-1) & MULT_106(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(48)<=signed(MULT_105(48)(MULT_SIZE-1) & MULT_105(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(48)(MULT_SIZE-1) & MULT_106(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(49)<=signed(MULT_105(49)(MULT_SIZE-1) & MULT_105(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(49)(MULT_SIZE-1) & MULT_106(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(50)<=signed(MULT_105(50)(MULT_SIZE-1) & MULT_105(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(50)(MULT_SIZE-1) & MULT_106(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(51)<=signed(MULT_105(51)(MULT_SIZE-1) & MULT_105(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(51)(MULT_SIZE-1) & MULT_106(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(52)<=signed(MULT_105(52)(MULT_SIZE-1) & MULT_105(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(52)(MULT_SIZE-1) & MULT_106(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(53)<=signed(MULT_105(53)(MULT_SIZE-1) & MULT_105(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(53)(MULT_SIZE-1) & MULT_106(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(54)<=signed(MULT_105(54)(MULT_SIZE-1) & MULT_105(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(54)(MULT_SIZE-1) & MULT_106(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(55)<=signed(MULT_105(55)(MULT_SIZE-1) & MULT_105(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(55)(MULT_SIZE-1) & MULT_106(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(56)<=signed(MULT_105(56)(MULT_SIZE-1) & MULT_105(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(56)(MULT_SIZE-1) & MULT_106(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(57)<=signed(MULT_105(57)(MULT_SIZE-1) & MULT_105(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(57)(MULT_SIZE-1) & MULT_106(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(58)<=signed(MULT_105(58)(MULT_SIZE-1) & MULT_105(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(58)(MULT_SIZE-1) & MULT_106(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(59)<=signed(MULT_105(59)(MULT_SIZE-1) & MULT_105(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(59)(MULT_SIZE-1) & MULT_106(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(60)<=signed(MULT_105(60)(MULT_SIZE-1) & MULT_105(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(60)(MULT_SIZE-1) & MULT_106(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(61)<=signed(MULT_105(61)(MULT_SIZE-1) & MULT_105(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(61)(MULT_SIZE-1) & MULT_106(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(62)<=signed(MULT_105(62)(MULT_SIZE-1) & MULT_105(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(62)(MULT_SIZE-1) & MULT_106(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(63)<=signed(MULT_105(63)(MULT_SIZE-1) & MULT_105(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(63)(MULT_SIZE-1) & MULT_106(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(64)<=signed(MULT_105(64)(MULT_SIZE-1) & MULT_105(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(64)(MULT_SIZE-1) & MULT_106(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(65)<=signed(MULT_105(65)(MULT_SIZE-1) & MULT_105(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(65)(MULT_SIZE-1) & MULT_106(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(66)<=signed(MULT_105(66)(MULT_SIZE-1) & MULT_105(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(66)(MULT_SIZE-1) & MULT_106(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(67)<=signed(MULT_105(67)(MULT_SIZE-1) & MULT_105(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(67)(MULT_SIZE-1) & MULT_106(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(68)<=signed(MULT_105(68)(MULT_SIZE-1) & MULT_105(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(68)(MULT_SIZE-1) & MULT_106(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(69)<=signed(MULT_105(69)(MULT_SIZE-1) & MULT_105(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(69)(MULT_SIZE-1) & MULT_106(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(70)<=signed(MULT_105(70)(MULT_SIZE-1) & MULT_105(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(70)(MULT_SIZE-1) & MULT_106(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(71)<=signed(MULT_105(71)(MULT_SIZE-1) & MULT_105(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(71)(MULT_SIZE-1) & MULT_106(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(72)<=signed(MULT_105(72)(MULT_SIZE-1) & MULT_105(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(72)(MULT_SIZE-1) & MULT_106(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(73)<=signed(MULT_105(73)(MULT_SIZE-1) & MULT_105(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(73)(MULT_SIZE-1) & MULT_106(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(74)<=signed(MULT_105(74)(MULT_SIZE-1) & MULT_105(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(74)(MULT_SIZE-1) & MULT_106(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(75)<=signed(MULT_105(75)(MULT_SIZE-1) & MULT_105(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(75)(MULT_SIZE-1) & MULT_106(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(76)<=signed(MULT_105(76)(MULT_SIZE-1) & MULT_105(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(76)(MULT_SIZE-1) & MULT_106(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(77)<=signed(MULT_105(77)(MULT_SIZE-1) & MULT_105(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(77)(MULT_SIZE-1) & MULT_106(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(78)<=signed(MULT_105(78)(MULT_SIZE-1) & MULT_105(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(78)(MULT_SIZE-1) & MULT_106(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(79)<=signed(MULT_105(79)(MULT_SIZE-1) & MULT_105(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(79)(MULT_SIZE-1) & MULT_106(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(80)<=signed(MULT_105(80)(MULT_SIZE-1) & MULT_105(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(80)(MULT_SIZE-1) & MULT_106(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(81)<=signed(MULT_105(81)(MULT_SIZE-1) & MULT_105(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(81)(MULT_SIZE-1) & MULT_106(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(82)<=signed(MULT_105(82)(MULT_SIZE-1) & MULT_105(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(82)(MULT_SIZE-1) & MULT_106(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_53(83)<=signed(MULT_105(83)(MULT_SIZE-1) & MULT_105(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_106(83)(MULT_SIZE-1) & MULT_106(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_54(0)<=signed(MULT_107(0)(MULT_SIZE-1) & MULT_107(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(0)(MULT_SIZE-1) & MULT_108(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(1)<=signed(MULT_107(1)(MULT_SIZE-1) & MULT_107(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(1)(MULT_SIZE-1) & MULT_108(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(2)<=signed(MULT_107(2)(MULT_SIZE-1) & MULT_107(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(2)(MULT_SIZE-1) & MULT_108(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(3)<=signed(MULT_107(3)(MULT_SIZE-1) & MULT_107(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(3)(MULT_SIZE-1) & MULT_108(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(4)<=signed(MULT_107(4)(MULT_SIZE-1) & MULT_107(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(4)(MULT_SIZE-1) & MULT_108(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(5)<=signed(MULT_107(5)(MULT_SIZE-1) & MULT_107(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(5)(MULT_SIZE-1) & MULT_108(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(6)<=signed(MULT_107(6)(MULT_SIZE-1) & MULT_107(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(6)(MULT_SIZE-1) & MULT_108(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(7)<=signed(MULT_107(7)(MULT_SIZE-1) & MULT_107(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(7)(MULT_SIZE-1) & MULT_108(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(8)<=signed(MULT_107(8)(MULT_SIZE-1) & MULT_107(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(8)(MULT_SIZE-1) & MULT_108(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(9)<=signed(MULT_107(9)(MULT_SIZE-1) & MULT_107(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(9)(MULT_SIZE-1) & MULT_108(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(10)<=signed(MULT_107(10)(MULT_SIZE-1) & MULT_107(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(10)(MULT_SIZE-1) & MULT_108(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(11)<=signed(MULT_107(11)(MULT_SIZE-1) & MULT_107(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(11)(MULT_SIZE-1) & MULT_108(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(12)<=signed(MULT_107(12)(MULT_SIZE-1) & MULT_107(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(12)(MULT_SIZE-1) & MULT_108(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(13)<=signed(MULT_107(13)(MULT_SIZE-1) & MULT_107(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(13)(MULT_SIZE-1) & MULT_108(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(14)<=signed(MULT_107(14)(MULT_SIZE-1) & MULT_107(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(14)(MULT_SIZE-1) & MULT_108(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(15)<=signed(MULT_107(15)(MULT_SIZE-1) & MULT_107(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(15)(MULT_SIZE-1) & MULT_108(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(16)<=signed(MULT_107(16)(MULT_SIZE-1) & MULT_107(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(16)(MULT_SIZE-1) & MULT_108(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(17)<=signed(MULT_107(17)(MULT_SIZE-1) & MULT_107(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(17)(MULT_SIZE-1) & MULT_108(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(18)<=signed(MULT_107(18)(MULT_SIZE-1) & MULT_107(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(18)(MULT_SIZE-1) & MULT_108(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(19)<=signed(MULT_107(19)(MULT_SIZE-1) & MULT_107(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(19)(MULT_SIZE-1) & MULT_108(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(20)<=signed(MULT_107(20)(MULT_SIZE-1) & MULT_107(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(20)(MULT_SIZE-1) & MULT_108(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(21)<=signed(MULT_107(21)(MULT_SIZE-1) & MULT_107(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(21)(MULT_SIZE-1) & MULT_108(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(22)<=signed(MULT_107(22)(MULT_SIZE-1) & MULT_107(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(22)(MULT_SIZE-1) & MULT_108(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(23)<=signed(MULT_107(23)(MULT_SIZE-1) & MULT_107(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(23)(MULT_SIZE-1) & MULT_108(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(24)<=signed(MULT_107(24)(MULT_SIZE-1) & MULT_107(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(24)(MULT_SIZE-1) & MULT_108(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(25)<=signed(MULT_107(25)(MULT_SIZE-1) & MULT_107(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(25)(MULT_SIZE-1) & MULT_108(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(26)<=signed(MULT_107(26)(MULT_SIZE-1) & MULT_107(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(26)(MULT_SIZE-1) & MULT_108(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(27)<=signed(MULT_107(27)(MULT_SIZE-1) & MULT_107(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(27)(MULT_SIZE-1) & MULT_108(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(28)<=signed(MULT_107(28)(MULT_SIZE-1) & MULT_107(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(28)(MULT_SIZE-1) & MULT_108(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(29)<=signed(MULT_107(29)(MULT_SIZE-1) & MULT_107(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(29)(MULT_SIZE-1) & MULT_108(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(30)<=signed(MULT_107(30)(MULT_SIZE-1) & MULT_107(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(30)(MULT_SIZE-1) & MULT_108(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(31)<=signed(MULT_107(31)(MULT_SIZE-1) & MULT_107(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(31)(MULT_SIZE-1) & MULT_108(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(32)<=signed(MULT_107(32)(MULT_SIZE-1) & MULT_107(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(32)(MULT_SIZE-1) & MULT_108(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(33)<=signed(MULT_107(33)(MULT_SIZE-1) & MULT_107(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(33)(MULT_SIZE-1) & MULT_108(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(34)<=signed(MULT_107(34)(MULT_SIZE-1) & MULT_107(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(34)(MULT_SIZE-1) & MULT_108(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(35)<=signed(MULT_107(35)(MULT_SIZE-1) & MULT_107(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(35)(MULT_SIZE-1) & MULT_108(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(36)<=signed(MULT_107(36)(MULT_SIZE-1) & MULT_107(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(36)(MULT_SIZE-1) & MULT_108(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(37)<=signed(MULT_107(37)(MULT_SIZE-1) & MULT_107(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(37)(MULT_SIZE-1) & MULT_108(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(38)<=signed(MULT_107(38)(MULT_SIZE-1) & MULT_107(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(38)(MULT_SIZE-1) & MULT_108(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(39)<=signed(MULT_107(39)(MULT_SIZE-1) & MULT_107(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(39)(MULT_SIZE-1) & MULT_108(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(40)<=signed(MULT_107(40)(MULT_SIZE-1) & MULT_107(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(40)(MULT_SIZE-1) & MULT_108(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(41)<=signed(MULT_107(41)(MULT_SIZE-1) & MULT_107(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(41)(MULT_SIZE-1) & MULT_108(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(42)<=signed(MULT_107(42)(MULT_SIZE-1) & MULT_107(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(42)(MULT_SIZE-1) & MULT_108(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(43)<=signed(MULT_107(43)(MULT_SIZE-1) & MULT_107(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(43)(MULT_SIZE-1) & MULT_108(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(44)<=signed(MULT_107(44)(MULT_SIZE-1) & MULT_107(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(44)(MULT_SIZE-1) & MULT_108(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(45)<=signed(MULT_107(45)(MULT_SIZE-1) & MULT_107(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(45)(MULT_SIZE-1) & MULT_108(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(46)<=signed(MULT_107(46)(MULT_SIZE-1) & MULT_107(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(46)(MULT_SIZE-1) & MULT_108(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(47)<=signed(MULT_107(47)(MULT_SIZE-1) & MULT_107(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(47)(MULT_SIZE-1) & MULT_108(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(48)<=signed(MULT_107(48)(MULT_SIZE-1) & MULT_107(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(48)(MULT_SIZE-1) & MULT_108(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(49)<=signed(MULT_107(49)(MULT_SIZE-1) & MULT_107(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(49)(MULT_SIZE-1) & MULT_108(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(50)<=signed(MULT_107(50)(MULT_SIZE-1) & MULT_107(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(50)(MULT_SIZE-1) & MULT_108(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(51)<=signed(MULT_107(51)(MULT_SIZE-1) & MULT_107(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(51)(MULT_SIZE-1) & MULT_108(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(52)<=signed(MULT_107(52)(MULT_SIZE-1) & MULT_107(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(52)(MULT_SIZE-1) & MULT_108(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(53)<=signed(MULT_107(53)(MULT_SIZE-1) & MULT_107(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(53)(MULT_SIZE-1) & MULT_108(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(54)<=signed(MULT_107(54)(MULT_SIZE-1) & MULT_107(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(54)(MULT_SIZE-1) & MULT_108(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(55)<=signed(MULT_107(55)(MULT_SIZE-1) & MULT_107(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(55)(MULT_SIZE-1) & MULT_108(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(56)<=signed(MULT_107(56)(MULT_SIZE-1) & MULT_107(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(56)(MULT_SIZE-1) & MULT_108(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(57)<=signed(MULT_107(57)(MULT_SIZE-1) & MULT_107(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(57)(MULT_SIZE-1) & MULT_108(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(58)<=signed(MULT_107(58)(MULT_SIZE-1) & MULT_107(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(58)(MULT_SIZE-1) & MULT_108(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(59)<=signed(MULT_107(59)(MULT_SIZE-1) & MULT_107(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(59)(MULT_SIZE-1) & MULT_108(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(60)<=signed(MULT_107(60)(MULT_SIZE-1) & MULT_107(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(60)(MULT_SIZE-1) & MULT_108(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(61)<=signed(MULT_107(61)(MULT_SIZE-1) & MULT_107(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(61)(MULT_SIZE-1) & MULT_108(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(62)<=signed(MULT_107(62)(MULT_SIZE-1) & MULT_107(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(62)(MULT_SIZE-1) & MULT_108(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(63)<=signed(MULT_107(63)(MULT_SIZE-1) & MULT_107(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(63)(MULT_SIZE-1) & MULT_108(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(64)<=signed(MULT_107(64)(MULT_SIZE-1) & MULT_107(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(64)(MULT_SIZE-1) & MULT_108(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(65)<=signed(MULT_107(65)(MULT_SIZE-1) & MULT_107(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(65)(MULT_SIZE-1) & MULT_108(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(66)<=signed(MULT_107(66)(MULT_SIZE-1) & MULT_107(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(66)(MULT_SIZE-1) & MULT_108(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(67)<=signed(MULT_107(67)(MULT_SIZE-1) & MULT_107(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(67)(MULT_SIZE-1) & MULT_108(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(68)<=signed(MULT_107(68)(MULT_SIZE-1) & MULT_107(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(68)(MULT_SIZE-1) & MULT_108(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(69)<=signed(MULT_107(69)(MULT_SIZE-1) & MULT_107(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(69)(MULT_SIZE-1) & MULT_108(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(70)<=signed(MULT_107(70)(MULT_SIZE-1) & MULT_107(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(70)(MULT_SIZE-1) & MULT_108(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(71)<=signed(MULT_107(71)(MULT_SIZE-1) & MULT_107(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(71)(MULT_SIZE-1) & MULT_108(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(72)<=signed(MULT_107(72)(MULT_SIZE-1) & MULT_107(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(72)(MULT_SIZE-1) & MULT_108(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(73)<=signed(MULT_107(73)(MULT_SIZE-1) & MULT_107(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(73)(MULT_SIZE-1) & MULT_108(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(74)<=signed(MULT_107(74)(MULT_SIZE-1) & MULT_107(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(74)(MULT_SIZE-1) & MULT_108(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(75)<=signed(MULT_107(75)(MULT_SIZE-1) & MULT_107(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(75)(MULT_SIZE-1) & MULT_108(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(76)<=signed(MULT_107(76)(MULT_SIZE-1) & MULT_107(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(76)(MULT_SIZE-1) & MULT_108(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(77)<=signed(MULT_107(77)(MULT_SIZE-1) & MULT_107(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(77)(MULT_SIZE-1) & MULT_108(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(78)<=signed(MULT_107(78)(MULT_SIZE-1) & MULT_107(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(78)(MULT_SIZE-1) & MULT_108(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(79)<=signed(MULT_107(79)(MULT_SIZE-1) & MULT_107(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(79)(MULT_SIZE-1) & MULT_108(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(80)<=signed(MULT_107(80)(MULT_SIZE-1) & MULT_107(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(80)(MULT_SIZE-1) & MULT_108(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(81)<=signed(MULT_107(81)(MULT_SIZE-1) & MULT_107(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(81)(MULT_SIZE-1) & MULT_108(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(82)<=signed(MULT_107(82)(MULT_SIZE-1) & MULT_107(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(82)(MULT_SIZE-1) & MULT_108(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_54(83)<=signed(MULT_107(83)(MULT_SIZE-1) & MULT_107(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_108(83)(MULT_SIZE-1) & MULT_108(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_55(0)<=signed(MULT_109(0)(MULT_SIZE-1) & MULT_109(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(0)(MULT_SIZE-1) & MULT_110(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(1)<=signed(MULT_109(1)(MULT_SIZE-1) & MULT_109(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(1)(MULT_SIZE-1) & MULT_110(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(2)<=signed(MULT_109(2)(MULT_SIZE-1) & MULT_109(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(2)(MULT_SIZE-1) & MULT_110(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(3)<=signed(MULT_109(3)(MULT_SIZE-1) & MULT_109(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(3)(MULT_SIZE-1) & MULT_110(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(4)<=signed(MULT_109(4)(MULT_SIZE-1) & MULT_109(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(4)(MULT_SIZE-1) & MULT_110(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(5)<=signed(MULT_109(5)(MULT_SIZE-1) & MULT_109(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(5)(MULT_SIZE-1) & MULT_110(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(6)<=signed(MULT_109(6)(MULT_SIZE-1) & MULT_109(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(6)(MULT_SIZE-1) & MULT_110(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(7)<=signed(MULT_109(7)(MULT_SIZE-1) & MULT_109(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(7)(MULT_SIZE-1) & MULT_110(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(8)<=signed(MULT_109(8)(MULT_SIZE-1) & MULT_109(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(8)(MULT_SIZE-1) & MULT_110(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(9)<=signed(MULT_109(9)(MULT_SIZE-1) & MULT_109(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(9)(MULT_SIZE-1) & MULT_110(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(10)<=signed(MULT_109(10)(MULT_SIZE-1) & MULT_109(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(10)(MULT_SIZE-1) & MULT_110(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(11)<=signed(MULT_109(11)(MULT_SIZE-1) & MULT_109(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(11)(MULT_SIZE-1) & MULT_110(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(12)<=signed(MULT_109(12)(MULT_SIZE-1) & MULT_109(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(12)(MULT_SIZE-1) & MULT_110(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(13)<=signed(MULT_109(13)(MULT_SIZE-1) & MULT_109(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(13)(MULT_SIZE-1) & MULT_110(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(14)<=signed(MULT_109(14)(MULT_SIZE-1) & MULT_109(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(14)(MULT_SIZE-1) & MULT_110(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(15)<=signed(MULT_109(15)(MULT_SIZE-1) & MULT_109(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(15)(MULT_SIZE-1) & MULT_110(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(16)<=signed(MULT_109(16)(MULT_SIZE-1) & MULT_109(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(16)(MULT_SIZE-1) & MULT_110(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(17)<=signed(MULT_109(17)(MULT_SIZE-1) & MULT_109(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(17)(MULT_SIZE-1) & MULT_110(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(18)<=signed(MULT_109(18)(MULT_SIZE-1) & MULT_109(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(18)(MULT_SIZE-1) & MULT_110(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(19)<=signed(MULT_109(19)(MULT_SIZE-1) & MULT_109(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(19)(MULT_SIZE-1) & MULT_110(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(20)<=signed(MULT_109(20)(MULT_SIZE-1) & MULT_109(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(20)(MULT_SIZE-1) & MULT_110(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(21)<=signed(MULT_109(21)(MULT_SIZE-1) & MULT_109(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(21)(MULT_SIZE-1) & MULT_110(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(22)<=signed(MULT_109(22)(MULT_SIZE-1) & MULT_109(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(22)(MULT_SIZE-1) & MULT_110(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(23)<=signed(MULT_109(23)(MULT_SIZE-1) & MULT_109(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(23)(MULT_SIZE-1) & MULT_110(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(24)<=signed(MULT_109(24)(MULT_SIZE-1) & MULT_109(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(24)(MULT_SIZE-1) & MULT_110(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(25)<=signed(MULT_109(25)(MULT_SIZE-1) & MULT_109(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(25)(MULT_SIZE-1) & MULT_110(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(26)<=signed(MULT_109(26)(MULT_SIZE-1) & MULT_109(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(26)(MULT_SIZE-1) & MULT_110(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(27)<=signed(MULT_109(27)(MULT_SIZE-1) & MULT_109(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(27)(MULT_SIZE-1) & MULT_110(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(28)<=signed(MULT_109(28)(MULT_SIZE-1) & MULT_109(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(28)(MULT_SIZE-1) & MULT_110(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(29)<=signed(MULT_109(29)(MULT_SIZE-1) & MULT_109(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(29)(MULT_SIZE-1) & MULT_110(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(30)<=signed(MULT_109(30)(MULT_SIZE-1) & MULT_109(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(30)(MULT_SIZE-1) & MULT_110(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(31)<=signed(MULT_109(31)(MULT_SIZE-1) & MULT_109(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(31)(MULT_SIZE-1) & MULT_110(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(32)<=signed(MULT_109(32)(MULT_SIZE-1) & MULT_109(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(32)(MULT_SIZE-1) & MULT_110(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(33)<=signed(MULT_109(33)(MULT_SIZE-1) & MULT_109(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(33)(MULT_SIZE-1) & MULT_110(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(34)<=signed(MULT_109(34)(MULT_SIZE-1) & MULT_109(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(34)(MULT_SIZE-1) & MULT_110(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(35)<=signed(MULT_109(35)(MULT_SIZE-1) & MULT_109(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(35)(MULT_SIZE-1) & MULT_110(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(36)<=signed(MULT_109(36)(MULT_SIZE-1) & MULT_109(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(36)(MULT_SIZE-1) & MULT_110(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(37)<=signed(MULT_109(37)(MULT_SIZE-1) & MULT_109(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(37)(MULT_SIZE-1) & MULT_110(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(38)<=signed(MULT_109(38)(MULT_SIZE-1) & MULT_109(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(38)(MULT_SIZE-1) & MULT_110(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(39)<=signed(MULT_109(39)(MULT_SIZE-1) & MULT_109(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(39)(MULT_SIZE-1) & MULT_110(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(40)<=signed(MULT_109(40)(MULT_SIZE-1) & MULT_109(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(40)(MULT_SIZE-1) & MULT_110(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(41)<=signed(MULT_109(41)(MULT_SIZE-1) & MULT_109(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(41)(MULT_SIZE-1) & MULT_110(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(42)<=signed(MULT_109(42)(MULT_SIZE-1) & MULT_109(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(42)(MULT_SIZE-1) & MULT_110(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(43)<=signed(MULT_109(43)(MULT_SIZE-1) & MULT_109(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(43)(MULT_SIZE-1) & MULT_110(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(44)<=signed(MULT_109(44)(MULT_SIZE-1) & MULT_109(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(44)(MULT_SIZE-1) & MULT_110(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(45)<=signed(MULT_109(45)(MULT_SIZE-1) & MULT_109(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(45)(MULT_SIZE-1) & MULT_110(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(46)<=signed(MULT_109(46)(MULT_SIZE-1) & MULT_109(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(46)(MULT_SIZE-1) & MULT_110(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(47)<=signed(MULT_109(47)(MULT_SIZE-1) & MULT_109(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(47)(MULT_SIZE-1) & MULT_110(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(48)<=signed(MULT_109(48)(MULT_SIZE-1) & MULT_109(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(48)(MULT_SIZE-1) & MULT_110(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(49)<=signed(MULT_109(49)(MULT_SIZE-1) & MULT_109(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(49)(MULT_SIZE-1) & MULT_110(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(50)<=signed(MULT_109(50)(MULT_SIZE-1) & MULT_109(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(50)(MULT_SIZE-1) & MULT_110(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(51)<=signed(MULT_109(51)(MULT_SIZE-1) & MULT_109(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(51)(MULT_SIZE-1) & MULT_110(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(52)<=signed(MULT_109(52)(MULT_SIZE-1) & MULT_109(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(52)(MULT_SIZE-1) & MULT_110(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(53)<=signed(MULT_109(53)(MULT_SIZE-1) & MULT_109(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(53)(MULT_SIZE-1) & MULT_110(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(54)<=signed(MULT_109(54)(MULT_SIZE-1) & MULT_109(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(54)(MULT_SIZE-1) & MULT_110(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(55)<=signed(MULT_109(55)(MULT_SIZE-1) & MULT_109(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(55)(MULT_SIZE-1) & MULT_110(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(56)<=signed(MULT_109(56)(MULT_SIZE-1) & MULT_109(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(56)(MULT_SIZE-1) & MULT_110(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(57)<=signed(MULT_109(57)(MULT_SIZE-1) & MULT_109(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(57)(MULT_SIZE-1) & MULT_110(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(58)<=signed(MULT_109(58)(MULT_SIZE-1) & MULT_109(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(58)(MULT_SIZE-1) & MULT_110(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(59)<=signed(MULT_109(59)(MULT_SIZE-1) & MULT_109(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(59)(MULT_SIZE-1) & MULT_110(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(60)<=signed(MULT_109(60)(MULT_SIZE-1) & MULT_109(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(60)(MULT_SIZE-1) & MULT_110(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(61)<=signed(MULT_109(61)(MULT_SIZE-1) & MULT_109(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(61)(MULT_SIZE-1) & MULT_110(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(62)<=signed(MULT_109(62)(MULT_SIZE-1) & MULT_109(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(62)(MULT_SIZE-1) & MULT_110(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(63)<=signed(MULT_109(63)(MULT_SIZE-1) & MULT_109(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(63)(MULT_SIZE-1) & MULT_110(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(64)<=signed(MULT_109(64)(MULT_SIZE-1) & MULT_109(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(64)(MULT_SIZE-1) & MULT_110(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(65)<=signed(MULT_109(65)(MULT_SIZE-1) & MULT_109(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(65)(MULT_SIZE-1) & MULT_110(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(66)<=signed(MULT_109(66)(MULT_SIZE-1) & MULT_109(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(66)(MULT_SIZE-1) & MULT_110(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(67)<=signed(MULT_109(67)(MULT_SIZE-1) & MULT_109(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(67)(MULT_SIZE-1) & MULT_110(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(68)<=signed(MULT_109(68)(MULT_SIZE-1) & MULT_109(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(68)(MULT_SIZE-1) & MULT_110(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(69)<=signed(MULT_109(69)(MULT_SIZE-1) & MULT_109(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(69)(MULT_SIZE-1) & MULT_110(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(70)<=signed(MULT_109(70)(MULT_SIZE-1) & MULT_109(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(70)(MULT_SIZE-1) & MULT_110(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(71)<=signed(MULT_109(71)(MULT_SIZE-1) & MULT_109(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(71)(MULT_SIZE-1) & MULT_110(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(72)<=signed(MULT_109(72)(MULT_SIZE-1) & MULT_109(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(72)(MULT_SIZE-1) & MULT_110(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(73)<=signed(MULT_109(73)(MULT_SIZE-1) & MULT_109(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(73)(MULT_SIZE-1) & MULT_110(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(74)<=signed(MULT_109(74)(MULT_SIZE-1) & MULT_109(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(74)(MULT_SIZE-1) & MULT_110(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(75)<=signed(MULT_109(75)(MULT_SIZE-1) & MULT_109(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(75)(MULT_SIZE-1) & MULT_110(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(76)<=signed(MULT_109(76)(MULT_SIZE-1) & MULT_109(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(76)(MULT_SIZE-1) & MULT_110(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(77)<=signed(MULT_109(77)(MULT_SIZE-1) & MULT_109(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(77)(MULT_SIZE-1) & MULT_110(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(78)<=signed(MULT_109(78)(MULT_SIZE-1) & MULT_109(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(78)(MULT_SIZE-1) & MULT_110(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(79)<=signed(MULT_109(79)(MULT_SIZE-1) & MULT_109(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(79)(MULT_SIZE-1) & MULT_110(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(80)<=signed(MULT_109(80)(MULT_SIZE-1) & MULT_109(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(80)(MULT_SIZE-1) & MULT_110(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(81)<=signed(MULT_109(81)(MULT_SIZE-1) & MULT_109(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(81)(MULT_SIZE-1) & MULT_110(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(82)<=signed(MULT_109(82)(MULT_SIZE-1) & MULT_109(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(82)(MULT_SIZE-1) & MULT_110(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_55(83)<=signed(MULT_109(83)(MULT_SIZE-1) & MULT_109(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_110(83)(MULT_SIZE-1) & MULT_110(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_56(0)<=signed(MULT_111(0)(MULT_SIZE-1) & MULT_111(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(0)(MULT_SIZE-1) & MULT_112(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(1)<=signed(MULT_111(1)(MULT_SIZE-1) & MULT_111(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(1)(MULT_SIZE-1) & MULT_112(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(2)<=signed(MULT_111(2)(MULT_SIZE-1) & MULT_111(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(2)(MULT_SIZE-1) & MULT_112(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(3)<=signed(MULT_111(3)(MULT_SIZE-1) & MULT_111(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(3)(MULT_SIZE-1) & MULT_112(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(4)<=signed(MULT_111(4)(MULT_SIZE-1) & MULT_111(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(4)(MULT_SIZE-1) & MULT_112(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(5)<=signed(MULT_111(5)(MULT_SIZE-1) & MULT_111(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(5)(MULT_SIZE-1) & MULT_112(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(6)<=signed(MULT_111(6)(MULT_SIZE-1) & MULT_111(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(6)(MULT_SIZE-1) & MULT_112(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(7)<=signed(MULT_111(7)(MULT_SIZE-1) & MULT_111(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(7)(MULT_SIZE-1) & MULT_112(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(8)<=signed(MULT_111(8)(MULT_SIZE-1) & MULT_111(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(8)(MULT_SIZE-1) & MULT_112(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(9)<=signed(MULT_111(9)(MULT_SIZE-1) & MULT_111(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(9)(MULT_SIZE-1) & MULT_112(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(10)<=signed(MULT_111(10)(MULT_SIZE-1) & MULT_111(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(10)(MULT_SIZE-1) & MULT_112(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(11)<=signed(MULT_111(11)(MULT_SIZE-1) & MULT_111(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(11)(MULT_SIZE-1) & MULT_112(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(12)<=signed(MULT_111(12)(MULT_SIZE-1) & MULT_111(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(12)(MULT_SIZE-1) & MULT_112(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(13)<=signed(MULT_111(13)(MULT_SIZE-1) & MULT_111(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(13)(MULT_SIZE-1) & MULT_112(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(14)<=signed(MULT_111(14)(MULT_SIZE-1) & MULT_111(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(14)(MULT_SIZE-1) & MULT_112(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(15)<=signed(MULT_111(15)(MULT_SIZE-1) & MULT_111(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(15)(MULT_SIZE-1) & MULT_112(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(16)<=signed(MULT_111(16)(MULT_SIZE-1) & MULT_111(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(16)(MULT_SIZE-1) & MULT_112(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(17)<=signed(MULT_111(17)(MULT_SIZE-1) & MULT_111(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(17)(MULT_SIZE-1) & MULT_112(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(18)<=signed(MULT_111(18)(MULT_SIZE-1) & MULT_111(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(18)(MULT_SIZE-1) & MULT_112(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(19)<=signed(MULT_111(19)(MULT_SIZE-1) & MULT_111(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(19)(MULT_SIZE-1) & MULT_112(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(20)<=signed(MULT_111(20)(MULT_SIZE-1) & MULT_111(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(20)(MULT_SIZE-1) & MULT_112(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(21)<=signed(MULT_111(21)(MULT_SIZE-1) & MULT_111(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(21)(MULT_SIZE-1) & MULT_112(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(22)<=signed(MULT_111(22)(MULT_SIZE-1) & MULT_111(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(22)(MULT_SIZE-1) & MULT_112(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(23)<=signed(MULT_111(23)(MULT_SIZE-1) & MULT_111(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(23)(MULT_SIZE-1) & MULT_112(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(24)<=signed(MULT_111(24)(MULT_SIZE-1) & MULT_111(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(24)(MULT_SIZE-1) & MULT_112(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(25)<=signed(MULT_111(25)(MULT_SIZE-1) & MULT_111(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(25)(MULT_SIZE-1) & MULT_112(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(26)<=signed(MULT_111(26)(MULT_SIZE-1) & MULT_111(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(26)(MULT_SIZE-1) & MULT_112(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(27)<=signed(MULT_111(27)(MULT_SIZE-1) & MULT_111(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(27)(MULT_SIZE-1) & MULT_112(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(28)<=signed(MULT_111(28)(MULT_SIZE-1) & MULT_111(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(28)(MULT_SIZE-1) & MULT_112(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(29)<=signed(MULT_111(29)(MULT_SIZE-1) & MULT_111(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(29)(MULT_SIZE-1) & MULT_112(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(30)<=signed(MULT_111(30)(MULT_SIZE-1) & MULT_111(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(30)(MULT_SIZE-1) & MULT_112(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(31)<=signed(MULT_111(31)(MULT_SIZE-1) & MULT_111(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(31)(MULT_SIZE-1) & MULT_112(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(32)<=signed(MULT_111(32)(MULT_SIZE-1) & MULT_111(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(32)(MULT_SIZE-1) & MULT_112(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(33)<=signed(MULT_111(33)(MULT_SIZE-1) & MULT_111(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(33)(MULT_SIZE-1) & MULT_112(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(34)<=signed(MULT_111(34)(MULT_SIZE-1) & MULT_111(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(34)(MULT_SIZE-1) & MULT_112(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(35)<=signed(MULT_111(35)(MULT_SIZE-1) & MULT_111(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(35)(MULT_SIZE-1) & MULT_112(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(36)<=signed(MULT_111(36)(MULT_SIZE-1) & MULT_111(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(36)(MULT_SIZE-1) & MULT_112(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(37)<=signed(MULT_111(37)(MULT_SIZE-1) & MULT_111(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(37)(MULT_SIZE-1) & MULT_112(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(38)<=signed(MULT_111(38)(MULT_SIZE-1) & MULT_111(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(38)(MULT_SIZE-1) & MULT_112(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(39)<=signed(MULT_111(39)(MULT_SIZE-1) & MULT_111(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(39)(MULT_SIZE-1) & MULT_112(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(40)<=signed(MULT_111(40)(MULT_SIZE-1) & MULT_111(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(40)(MULT_SIZE-1) & MULT_112(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(41)<=signed(MULT_111(41)(MULT_SIZE-1) & MULT_111(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(41)(MULT_SIZE-1) & MULT_112(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(42)<=signed(MULT_111(42)(MULT_SIZE-1) & MULT_111(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(42)(MULT_SIZE-1) & MULT_112(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(43)<=signed(MULT_111(43)(MULT_SIZE-1) & MULT_111(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(43)(MULT_SIZE-1) & MULT_112(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(44)<=signed(MULT_111(44)(MULT_SIZE-1) & MULT_111(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(44)(MULT_SIZE-1) & MULT_112(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(45)<=signed(MULT_111(45)(MULT_SIZE-1) & MULT_111(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(45)(MULT_SIZE-1) & MULT_112(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(46)<=signed(MULT_111(46)(MULT_SIZE-1) & MULT_111(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(46)(MULT_SIZE-1) & MULT_112(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(47)<=signed(MULT_111(47)(MULT_SIZE-1) & MULT_111(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(47)(MULT_SIZE-1) & MULT_112(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(48)<=signed(MULT_111(48)(MULT_SIZE-1) & MULT_111(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(48)(MULT_SIZE-1) & MULT_112(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(49)<=signed(MULT_111(49)(MULT_SIZE-1) & MULT_111(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(49)(MULT_SIZE-1) & MULT_112(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(50)<=signed(MULT_111(50)(MULT_SIZE-1) & MULT_111(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(50)(MULT_SIZE-1) & MULT_112(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(51)<=signed(MULT_111(51)(MULT_SIZE-1) & MULT_111(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(51)(MULT_SIZE-1) & MULT_112(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(52)<=signed(MULT_111(52)(MULT_SIZE-1) & MULT_111(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(52)(MULT_SIZE-1) & MULT_112(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(53)<=signed(MULT_111(53)(MULT_SIZE-1) & MULT_111(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(53)(MULT_SIZE-1) & MULT_112(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(54)<=signed(MULT_111(54)(MULT_SIZE-1) & MULT_111(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(54)(MULT_SIZE-1) & MULT_112(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(55)<=signed(MULT_111(55)(MULT_SIZE-1) & MULT_111(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(55)(MULT_SIZE-1) & MULT_112(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(56)<=signed(MULT_111(56)(MULT_SIZE-1) & MULT_111(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(56)(MULT_SIZE-1) & MULT_112(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(57)<=signed(MULT_111(57)(MULT_SIZE-1) & MULT_111(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(57)(MULT_SIZE-1) & MULT_112(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(58)<=signed(MULT_111(58)(MULT_SIZE-1) & MULT_111(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(58)(MULT_SIZE-1) & MULT_112(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(59)<=signed(MULT_111(59)(MULT_SIZE-1) & MULT_111(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(59)(MULT_SIZE-1) & MULT_112(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(60)<=signed(MULT_111(60)(MULT_SIZE-1) & MULT_111(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(60)(MULT_SIZE-1) & MULT_112(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(61)<=signed(MULT_111(61)(MULT_SIZE-1) & MULT_111(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(61)(MULT_SIZE-1) & MULT_112(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(62)<=signed(MULT_111(62)(MULT_SIZE-1) & MULT_111(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(62)(MULT_SIZE-1) & MULT_112(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(63)<=signed(MULT_111(63)(MULT_SIZE-1) & MULT_111(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(63)(MULT_SIZE-1) & MULT_112(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(64)<=signed(MULT_111(64)(MULT_SIZE-1) & MULT_111(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(64)(MULT_SIZE-1) & MULT_112(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(65)<=signed(MULT_111(65)(MULT_SIZE-1) & MULT_111(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(65)(MULT_SIZE-1) & MULT_112(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(66)<=signed(MULT_111(66)(MULT_SIZE-1) & MULT_111(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(66)(MULT_SIZE-1) & MULT_112(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(67)<=signed(MULT_111(67)(MULT_SIZE-1) & MULT_111(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(67)(MULT_SIZE-1) & MULT_112(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(68)<=signed(MULT_111(68)(MULT_SIZE-1) & MULT_111(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(68)(MULT_SIZE-1) & MULT_112(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(69)<=signed(MULT_111(69)(MULT_SIZE-1) & MULT_111(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(69)(MULT_SIZE-1) & MULT_112(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(70)<=signed(MULT_111(70)(MULT_SIZE-1) & MULT_111(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(70)(MULT_SIZE-1) & MULT_112(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(71)<=signed(MULT_111(71)(MULT_SIZE-1) & MULT_111(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(71)(MULT_SIZE-1) & MULT_112(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(72)<=signed(MULT_111(72)(MULT_SIZE-1) & MULT_111(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(72)(MULT_SIZE-1) & MULT_112(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(73)<=signed(MULT_111(73)(MULT_SIZE-1) & MULT_111(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(73)(MULT_SIZE-1) & MULT_112(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(74)<=signed(MULT_111(74)(MULT_SIZE-1) & MULT_111(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(74)(MULT_SIZE-1) & MULT_112(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(75)<=signed(MULT_111(75)(MULT_SIZE-1) & MULT_111(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(75)(MULT_SIZE-1) & MULT_112(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(76)<=signed(MULT_111(76)(MULT_SIZE-1) & MULT_111(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(76)(MULT_SIZE-1) & MULT_112(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(77)<=signed(MULT_111(77)(MULT_SIZE-1) & MULT_111(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(77)(MULT_SIZE-1) & MULT_112(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(78)<=signed(MULT_111(78)(MULT_SIZE-1) & MULT_111(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(78)(MULT_SIZE-1) & MULT_112(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(79)<=signed(MULT_111(79)(MULT_SIZE-1) & MULT_111(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(79)(MULT_SIZE-1) & MULT_112(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(80)<=signed(MULT_111(80)(MULT_SIZE-1) & MULT_111(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(80)(MULT_SIZE-1) & MULT_112(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(81)<=signed(MULT_111(81)(MULT_SIZE-1) & MULT_111(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(81)(MULT_SIZE-1) & MULT_112(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(82)<=signed(MULT_111(82)(MULT_SIZE-1) & MULT_111(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(82)(MULT_SIZE-1) & MULT_112(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_56(83)<=signed(MULT_111(83)(MULT_SIZE-1) & MULT_111(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_112(83)(MULT_SIZE-1) & MULT_112(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_57(0)<=signed(MULT_113(0)(MULT_SIZE-1) & MULT_113(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(0)(MULT_SIZE-1) & MULT_114(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(1)<=signed(MULT_113(1)(MULT_SIZE-1) & MULT_113(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(1)(MULT_SIZE-1) & MULT_114(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(2)<=signed(MULT_113(2)(MULT_SIZE-1) & MULT_113(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(2)(MULT_SIZE-1) & MULT_114(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(3)<=signed(MULT_113(3)(MULT_SIZE-1) & MULT_113(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(3)(MULT_SIZE-1) & MULT_114(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(4)<=signed(MULT_113(4)(MULT_SIZE-1) & MULT_113(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(4)(MULT_SIZE-1) & MULT_114(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(5)<=signed(MULT_113(5)(MULT_SIZE-1) & MULT_113(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(5)(MULT_SIZE-1) & MULT_114(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(6)<=signed(MULT_113(6)(MULT_SIZE-1) & MULT_113(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(6)(MULT_SIZE-1) & MULT_114(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(7)<=signed(MULT_113(7)(MULT_SIZE-1) & MULT_113(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(7)(MULT_SIZE-1) & MULT_114(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(8)<=signed(MULT_113(8)(MULT_SIZE-1) & MULT_113(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(8)(MULT_SIZE-1) & MULT_114(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(9)<=signed(MULT_113(9)(MULT_SIZE-1) & MULT_113(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(9)(MULT_SIZE-1) & MULT_114(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(10)<=signed(MULT_113(10)(MULT_SIZE-1) & MULT_113(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(10)(MULT_SIZE-1) & MULT_114(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(11)<=signed(MULT_113(11)(MULT_SIZE-1) & MULT_113(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(11)(MULT_SIZE-1) & MULT_114(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(12)<=signed(MULT_113(12)(MULT_SIZE-1) & MULT_113(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(12)(MULT_SIZE-1) & MULT_114(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(13)<=signed(MULT_113(13)(MULT_SIZE-1) & MULT_113(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(13)(MULT_SIZE-1) & MULT_114(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(14)<=signed(MULT_113(14)(MULT_SIZE-1) & MULT_113(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(14)(MULT_SIZE-1) & MULT_114(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(15)<=signed(MULT_113(15)(MULT_SIZE-1) & MULT_113(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(15)(MULT_SIZE-1) & MULT_114(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(16)<=signed(MULT_113(16)(MULT_SIZE-1) & MULT_113(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(16)(MULT_SIZE-1) & MULT_114(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(17)<=signed(MULT_113(17)(MULT_SIZE-1) & MULT_113(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(17)(MULT_SIZE-1) & MULT_114(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(18)<=signed(MULT_113(18)(MULT_SIZE-1) & MULT_113(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(18)(MULT_SIZE-1) & MULT_114(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(19)<=signed(MULT_113(19)(MULT_SIZE-1) & MULT_113(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(19)(MULT_SIZE-1) & MULT_114(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(20)<=signed(MULT_113(20)(MULT_SIZE-1) & MULT_113(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(20)(MULT_SIZE-1) & MULT_114(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(21)<=signed(MULT_113(21)(MULT_SIZE-1) & MULT_113(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(21)(MULT_SIZE-1) & MULT_114(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(22)<=signed(MULT_113(22)(MULT_SIZE-1) & MULT_113(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(22)(MULT_SIZE-1) & MULT_114(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(23)<=signed(MULT_113(23)(MULT_SIZE-1) & MULT_113(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(23)(MULT_SIZE-1) & MULT_114(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(24)<=signed(MULT_113(24)(MULT_SIZE-1) & MULT_113(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(24)(MULT_SIZE-1) & MULT_114(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(25)<=signed(MULT_113(25)(MULT_SIZE-1) & MULT_113(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(25)(MULT_SIZE-1) & MULT_114(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(26)<=signed(MULT_113(26)(MULT_SIZE-1) & MULT_113(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(26)(MULT_SIZE-1) & MULT_114(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(27)<=signed(MULT_113(27)(MULT_SIZE-1) & MULT_113(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(27)(MULT_SIZE-1) & MULT_114(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(28)<=signed(MULT_113(28)(MULT_SIZE-1) & MULT_113(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(28)(MULT_SIZE-1) & MULT_114(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(29)<=signed(MULT_113(29)(MULT_SIZE-1) & MULT_113(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(29)(MULT_SIZE-1) & MULT_114(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(30)<=signed(MULT_113(30)(MULT_SIZE-1) & MULT_113(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(30)(MULT_SIZE-1) & MULT_114(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(31)<=signed(MULT_113(31)(MULT_SIZE-1) & MULT_113(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(31)(MULT_SIZE-1) & MULT_114(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(32)<=signed(MULT_113(32)(MULT_SIZE-1) & MULT_113(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(32)(MULT_SIZE-1) & MULT_114(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(33)<=signed(MULT_113(33)(MULT_SIZE-1) & MULT_113(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(33)(MULT_SIZE-1) & MULT_114(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(34)<=signed(MULT_113(34)(MULT_SIZE-1) & MULT_113(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(34)(MULT_SIZE-1) & MULT_114(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(35)<=signed(MULT_113(35)(MULT_SIZE-1) & MULT_113(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(35)(MULT_SIZE-1) & MULT_114(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(36)<=signed(MULT_113(36)(MULT_SIZE-1) & MULT_113(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(36)(MULT_SIZE-1) & MULT_114(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(37)<=signed(MULT_113(37)(MULT_SIZE-1) & MULT_113(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(37)(MULT_SIZE-1) & MULT_114(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(38)<=signed(MULT_113(38)(MULT_SIZE-1) & MULT_113(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(38)(MULT_SIZE-1) & MULT_114(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(39)<=signed(MULT_113(39)(MULT_SIZE-1) & MULT_113(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(39)(MULT_SIZE-1) & MULT_114(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(40)<=signed(MULT_113(40)(MULT_SIZE-1) & MULT_113(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(40)(MULT_SIZE-1) & MULT_114(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(41)<=signed(MULT_113(41)(MULT_SIZE-1) & MULT_113(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(41)(MULT_SIZE-1) & MULT_114(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(42)<=signed(MULT_113(42)(MULT_SIZE-1) & MULT_113(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(42)(MULT_SIZE-1) & MULT_114(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(43)<=signed(MULT_113(43)(MULT_SIZE-1) & MULT_113(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(43)(MULT_SIZE-1) & MULT_114(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(44)<=signed(MULT_113(44)(MULT_SIZE-1) & MULT_113(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(44)(MULT_SIZE-1) & MULT_114(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(45)<=signed(MULT_113(45)(MULT_SIZE-1) & MULT_113(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(45)(MULT_SIZE-1) & MULT_114(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(46)<=signed(MULT_113(46)(MULT_SIZE-1) & MULT_113(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(46)(MULT_SIZE-1) & MULT_114(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(47)<=signed(MULT_113(47)(MULT_SIZE-1) & MULT_113(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(47)(MULT_SIZE-1) & MULT_114(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(48)<=signed(MULT_113(48)(MULT_SIZE-1) & MULT_113(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(48)(MULT_SIZE-1) & MULT_114(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(49)<=signed(MULT_113(49)(MULT_SIZE-1) & MULT_113(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(49)(MULT_SIZE-1) & MULT_114(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(50)<=signed(MULT_113(50)(MULT_SIZE-1) & MULT_113(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(50)(MULT_SIZE-1) & MULT_114(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(51)<=signed(MULT_113(51)(MULT_SIZE-1) & MULT_113(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(51)(MULT_SIZE-1) & MULT_114(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(52)<=signed(MULT_113(52)(MULT_SIZE-1) & MULT_113(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(52)(MULT_SIZE-1) & MULT_114(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(53)<=signed(MULT_113(53)(MULT_SIZE-1) & MULT_113(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(53)(MULT_SIZE-1) & MULT_114(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(54)<=signed(MULT_113(54)(MULT_SIZE-1) & MULT_113(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(54)(MULT_SIZE-1) & MULT_114(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(55)<=signed(MULT_113(55)(MULT_SIZE-1) & MULT_113(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(55)(MULT_SIZE-1) & MULT_114(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(56)<=signed(MULT_113(56)(MULT_SIZE-1) & MULT_113(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(56)(MULT_SIZE-1) & MULT_114(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(57)<=signed(MULT_113(57)(MULT_SIZE-1) & MULT_113(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(57)(MULT_SIZE-1) & MULT_114(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(58)<=signed(MULT_113(58)(MULT_SIZE-1) & MULT_113(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(58)(MULT_SIZE-1) & MULT_114(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(59)<=signed(MULT_113(59)(MULT_SIZE-1) & MULT_113(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(59)(MULT_SIZE-1) & MULT_114(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(60)<=signed(MULT_113(60)(MULT_SIZE-1) & MULT_113(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(60)(MULT_SIZE-1) & MULT_114(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(61)<=signed(MULT_113(61)(MULT_SIZE-1) & MULT_113(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(61)(MULT_SIZE-1) & MULT_114(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(62)<=signed(MULT_113(62)(MULT_SIZE-1) & MULT_113(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(62)(MULT_SIZE-1) & MULT_114(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(63)<=signed(MULT_113(63)(MULT_SIZE-1) & MULT_113(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(63)(MULT_SIZE-1) & MULT_114(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(64)<=signed(MULT_113(64)(MULT_SIZE-1) & MULT_113(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(64)(MULT_SIZE-1) & MULT_114(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(65)<=signed(MULT_113(65)(MULT_SIZE-1) & MULT_113(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(65)(MULT_SIZE-1) & MULT_114(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(66)<=signed(MULT_113(66)(MULT_SIZE-1) & MULT_113(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(66)(MULT_SIZE-1) & MULT_114(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(67)<=signed(MULT_113(67)(MULT_SIZE-1) & MULT_113(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(67)(MULT_SIZE-1) & MULT_114(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(68)<=signed(MULT_113(68)(MULT_SIZE-1) & MULT_113(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(68)(MULT_SIZE-1) & MULT_114(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(69)<=signed(MULT_113(69)(MULT_SIZE-1) & MULT_113(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(69)(MULT_SIZE-1) & MULT_114(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(70)<=signed(MULT_113(70)(MULT_SIZE-1) & MULT_113(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(70)(MULT_SIZE-1) & MULT_114(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(71)<=signed(MULT_113(71)(MULT_SIZE-1) & MULT_113(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(71)(MULT_SIZE-1) & MULT_114(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(72)<=signed(MULT_113(72)(MULT_SIZE-1) & MULT_113(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(72)(MULT_SIZE-1) & MULT_114(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(73)<=signed(MULT_113(73)(MULT_SIZE-1) & MULT_113(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(73)(MULT_SIZE-1) & MULT_114(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(74)<=signed(MULT_113(74)(MULT_SIZE-1) & MULT_113(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(74)(MULT_SIZE-1) & MULT_114(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(75)<=signed(MULT_113(75)(MULT_SIZE-1) & MULT_113(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(75)(MULT_SIZE-1) & MULT_114(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(76)<=signed(MULT_113(76)(MULT_SIZE-1) & MULT_113(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(76)(MULT_SIZE-1) & MULT_114(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(77)<=signed(MULT_113(77)(MULT_SIZE-1) & MULT_113(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(77)(MULT_SIZE-1) & MULT_114(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(78)<=signed(MULT_113(78)(MULT_SIZE-1) & MULT_113(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(78)(MULT_SIZE-1) & MULT_114(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(79)<=signed(MULT_113(79)(MULT_SIZE-1) & MULT_113(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(79)(MULT_SIZE-1) & MULT_114(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(80)<=signed(MULT_113(80)(MULT_SIZE-1) & MULT_113(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(80)(MULT_SIZE-1) & MULT_114(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(81)<=signed(MULT_113(81)(MULT_SIZE-1) & MULT_113(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(81)(MULT_SIZE-1) & MULT_114(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(82)<=signed(MULT_113(82)(MULT_SIZE-1) & MULT_113(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(82)(MULT_SIZE-1) & MULT_114(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_57(83)<=signed(MULT_113(83)(MULT_SIZE-1) & MULT_113(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_114(83)(MULT_SIZE-1) & MULT_114(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_58(0)<=signed(MULT_115(0)(MULT_SIZE-1) & MULT_115(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(0)(MULT_SIZE-1) & MULT_116(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(1)<=signed(MULT_115(1)(MULT_SIZE-1) & MULT_115(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(1)(MULT_SIZE-1) & MULT_116(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(2)<=signed(MULT_115(2)(MULT_SIZE-1) & MULT_115(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(2)(MULT_SIZE-1) & MULT_116(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(3)<=signed(MULT_115(3)(MULT_SIZE-1) & MULT_115(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(3)(MULT_SIZE-1) & MULT_116(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(4)<=signed(MULT_115(4)(MULT_SIZE-1) & MULT_115(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(4)(MULT_SIZE-1) & MULT_116(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(5)<=signed(MULT_115(5)(MULT_SIZE-1) & MULT_115(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(5)(MULT_SIZE-1) & MULT_116(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(6)<=signed(MULT_115(6)(MULT_SIZE-1) & MULT_115(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(6)(MULT_SIZE-1) & MULT_116(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(7)<=signed(MULT_115(7)(MULT_SIZE-1) & MULT_115(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(7)(MULT_SIZE-1) & MULT_116(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(8)<=signed(MULT_115(8)(MULT_SIZE-1) & MULT_115(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(8)(MULT_SIZE-1) & MULT_116(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(9)<=signed(MULT_115(9)(MULT_SIZE-1) & MULT_115(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(9)(MULT_SIZE-1) & MULT_116(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(10)<=signed(MULT_115(10)(MULT_SIZE-1) & MULT_115(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(10)(MULT_SIZE-1) & MULT_116(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(11)<=signed(MULT_115(11)(MULT_SIZE-1) & MULT_115(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(11)(MULT_SIZE-1) & MULT_116(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(12)<=signed(MULT_115(12)(MULT_SIZE-1) & MULT_115(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(12)(MULT_SIZE-1) & MULT_116(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(13)<=signed(MULT_115(13)(MULT_SIZE-1) & MULT_115(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(13)(MULT_SIZE-1) & MULT_116(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(14)<=signed(MULT_115(14)(MULT_SIZE-1) & MULT_115(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(14)(MULT_SIZE-1) & MULT_116(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(15)<=signed(MULT_115(15)(MULT_SIZE-1) & MULT_115(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(15)(MULT_SIZE-1) & MULT_116(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(16)<=signed(MULT_115(16)(MULT_SIZE-1) & MULT_115(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(16)(MULT_SIZE-1) & MULT_116(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(17)<=signed(MULT_115(17)(MULT_SIZE-1) & MULT_115(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(17)(MULT_SIZE-1) & MULT_116(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(18)<=signed(MULT_115(18)(MULT_SIZE-1) & MULT_115(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(18)(MULT_SIZE-1) & MULT_116(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(19)<=signed(MULT_115(19)(MULT_SIZE-1) & MULT_115(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(19)(MULT_SIZE-1) & MULT_116(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(20)<=signed(MULT_115(20)(MULT_SIZE-1) & MULT_115(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(20)(MULT_SIZE-1) & MULT_116(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(21)<=signed(MULT_115(21)(MULT_SIZE-1) & MULT_115(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(21)(MULT_SIZE-1) & MULT_116(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(22)<=signed(MULT_115(22)(MULT_SIZE-1) & MULT_115(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(22)(MULT_SIZE-1) & MULT_116(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(23)<=signed(MULT_115(23)(MULT_SIZE-1) & MULT_115(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(23)(MULT_SIZE-1) & MULT_116(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(24)<=signed(MULT_115(24)(MULT_SIZE-1) & MULT_115(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(24)(MULT_SIZE-1) & MULT_116(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(25)<=signed(MULT_115(25)(MULT_SIZE-1) & MULT_115(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(25)(MULT_SIZE-1) & MULT_116(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(26)<=signed(MULT_115(26)(MULT_SIZE-1) & MULT_115(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(26)(MULT_SIZE-1) & MULT_116(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(27)<=signed(MULT_115(27)(MULT_SIZE-1) & MULT_115(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(27)(MULT_SIZE-1) & MULT_116(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(28)<=signed(MULT_115(28)(MULT_SIZE-1) & MULT_115(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(28)(MULT_SIZE-1) & MULT_116(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(29)<=signed(MULT_115(29)(MULT_SIZE-1) & MULT_115(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(29)(MULT_SIZE-1) & MULT_116(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(30)<=signed(MULT_115(30)(MULT_SIZE-1) & MULT_115(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(30)(MULT_SIZE-1) & MULT_116(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(31)<=signed(MULT_115(31)(MULT_SIZE-1) & MULT_115(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(31)(MULT_SIZE-1) & MULT_116(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(32)<=signed(MULT_115(32)(MULT_SIZE-1) & MULT_115(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(32)(MULT_SIZE-1) & MULT_116(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(33)<=signed(MULT_115(33)(MULT_SIZE-1) & MULT_115(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(33)(MULT_SIZE-1) & MULT_116(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(34)<=signed(MULT_115(34)(MULT_SIZE-1) & MULT_115(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(34)(MULT_SIZE-1) & MULT_116(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(35)<=signed(MULT_115(35)(MULT_SIZE-1) & MULT_115(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(35)(MULT_SIZE-1) & MULT_116(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(36)<=signed(MULT_115(36)(MULT_SIZE-1) & MULT_115(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(36)(MULT_SIZE-1) & MULT_116(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(37)<=signed(MULT_115(37)(MULT_SIZE-1) & MULT_115(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(37)(MULT_SIZE-1) & MULT_116(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(38)<=signed(MULT_115(38)(MULT_SIZE-1) & MULT_115(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(38)(MULT_SIZE-1) & MULT_116(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(39)<=signed(MULT_115(39)(MULT_SIZE-1) & MULT_115(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(39)(MULT_SIZE-1) & MULT_116(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(40)<=signed(MULT_115(40)(MULT_SIZE-1) & MULT_115(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(40)(MULT_SIZE-1) & MULT_116(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(41)<=signed(MULT_115(41)(MULT_SIZE-1) & MULT_115(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(41)(MULT_SIZE-1) & MULT_116(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(42)<=signed(MULT_115(42)(MULT_SIZE-1) & MULT_115(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(42)(MULT_SIZE-1) & MULT_116(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(43)<=signed(MULT_115(43)(MULT_SIZE-1) & MULT_115(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(43)(MULT_SIZE-1) & MULT_116(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(44)<=signed(MULT_115(44)(MULT_SIZE-1) & MULT_115(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(44)(MULT_SIZE-1) & MULT_116(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(45)<=signed(MULT_115(45)(MULT_SIZE-1) & MULT_115(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(45)(MULT_SIZE-1) & MULT_116(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(46)<=signed(MULT_115(46)(MULT_SIZE-1) & MULT_115(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(46)(MULT_SIZE-1) & MULT_116(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(47)<=signed(MULT_115(47)(MULT_SIZE-1) & MULT_115(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(47)(MULT_SIZE-1) & MULT_116(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(48)<=signed(MULT_115(48)(MULT_SIZE-1) & MULT_115(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(48)(MULT_SIZE-1) & MULT_116(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(49)<=signed(MULT_115(49)(MULT_SIZE-1) & MULT_115(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(49)(MULT_SIZE-1) & MULT_116(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(50)<=signed(MULT_115(50)(MULT_SIZE-1) & MULT_115(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(50)(MULT_SIZE-1) & MULT_116(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(51)<=signed(MULT_115(51)(MULT_SIZE-1) & MULT_115(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(51)(MULT_SIZE-1) & MULT_116(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(52)<=signed(MULT_115(52)(MULT_SIZE-1) & MULT_115(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(52)(MULT_SIZE-1) & MULT_116(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(53)<=signed(MULT_115(53)(MULT_SIZE-1) & MULT_115(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(53)(MULT_SIZE-1) & MULT_116(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(54)<=signed(MULT_115(54)(MULT_SIZE-1) & MULT_115(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(54)(MULT_SIZE-1) & MULT_116(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(55)<=signed(MULT_115(55)(MULT_SIZE-1) & MULT_115(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(55)(MULT_SIZE-1) & MULT_116(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(56)<=signed(MULT_115(56)(MULT_SIZE-1) & MULT_115(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(56)(MULT_SIZE-1) & MULT_116(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(57)<=signed(MULT_115(57)(MULT_SIZE-1) & MULT_115(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(57)(MULT_SIZE-1) & MULT_116(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(58)<=signed(MULT_115(58)(MULT_SIZE-1) & MULT_115(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(58)(MULT_SIZE-1) & MULT_116(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(59)<=signed(MULT_115(59)(MULT_SIZE-1) & MULT_115(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(59)(MULT_SIZE-1) & MULT_116(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(60)<=signed(MULT_115(60)(MULT_SIZE-1) & MULT_115(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(60)(MULT_SIZE-1) & MULT_116(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(61)<=signed(MULT_115(61)(MULT_SIZE-1) & MULT_115(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(61)(MULT_SIZE-1) & MULT_116(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(62)<=signed(MULT_115(62)(MULT_SIZE-1) & MULT_115(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(62)(MULT_SIZE-1) & MULT_116(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(63)<=signed(MULT_115(63)(MULT_SIZE-1) & MULT_115(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(63)(MULT_SIZE-1) & MULT_116(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(64)<=signed(MULT_115(64)(MULT_SIZE-1) & MULT_115(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(64)(MULT_SIZE-1) & MULT_116(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(65)<=signed(MULT_115(65)(MULT_SIZE-1) & MULT_115(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(65)(MULT_SIZE-1) & MULT_116(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(66)<=signed(MULT_115(66)(MULT_SIZE-1) & MULT_115(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(66)(MULT_SIZE-1) & MULT_116(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(67)<=signed(MULT_115(67)(MULT_SIZE-1) & MULT_115(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(67)(MULT_SIZE-1) & MULT_116(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(68)<=signed(MULT_115(68)(MULT_SIZE-1) & MULT_115(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(68)(MULT_SIZE-1) & MULT_116(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(69)<=signed(MULT_115(69)(MULT_SIZE-1) & MULT_115(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(69)(MULT_SIZE-1) & MULT_116(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(70)<=signed(MULT_115(70)(MULT_SIZE-1) & MULT_115(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(70)(MULT_SIZE-1) & MULT_116(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(71)<=signed(MULT_115(71)(MULT_SIZE-1) & MULT_115(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(71)(MULT_SIZE-1) & MULT_116(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(72)<=signed(MULT_115(72)(MULT_SIZE-1) & MULT_115(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(72)(MULT_SIZE-1) & MULT_116(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(73)<=signed(MULT_115(73)(MULT_SIZE-1) & MULT_115(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(73)(MULT_SIZE-1) & MULT_116(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(74)<=signed(MULT_115(74)(MULT_SIZE-1) & MULT_115(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(74)(MULT_SIZE-1) & MULT_116(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(75)<=signed(MULT_115(75)(MULT_SIZE-1) & MULT_115(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(75)(MULT_SIZE-1) & MULT_116(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(76)<=signed(MULT_115(76)(MULT_SIZE-1) & MULT_115(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(76)(MULT_SIZE-1) & MULT_116(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(77)<=signed(MULT_115(77)(MULT_SIZE-1) & MULT_115(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(77)(MULT_SIZE-1) & MULT_116(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(78)<=signed(MULT_115(78)(MULT_SIZE-1) & MULT_115(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(78)(MULT_SIZE-1) & MULT_116(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(79)<=signed(MULT_115(79)(MULT_SIZE-1) & MULT_115(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(79)(MULT_SIZE-1) & MULT_116(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(80)<=signed(MULT_115(80)(MULT_SIZE-1) & MULT_115(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(80)(MULT_SIZE-1) & MULT_116(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(81)<=signed(MULT_115(81)(MULT_SIZE-1) & MULT_115(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(81)(MULT_SIZE-1) & MULT_116(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(82)<=signed(MULT_115(82)(MULT_SIZE-1) & MULT_115(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(82)(MULT_SIZE-1) & MULT_116(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_58(83)<=signed(MULT_115(83)(MULT_SIZE-1) & MULT_115(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_116(83)(MULT_SIZE-1) & MULT_116(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_59(0)<=signed(MULT_117(0)(MULT_SIZE-1) & MULT_117(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(0)(MULT_SIZE-1) & MULT_118(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(1)<=signed(MULT_117(1)(MULT_SIZE-1) & MULT_117(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(1)(MULT_SIZE-1) & MULT_118(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(2)<=signed(MULT_117(2)(MULT_SIZE-1) & MULT_117(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(2)(MULT_SIZE-1) & MULT_118(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(3)<=signed(MULT_117(3)(MULT_SIZE-1) & MULT_117(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(3)(MULT_SIZE-1) & MULT_118(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(4)<=signed(MULT_117(4)(MULT_SIZE-1) & MULT_117(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(4)(MULT_SIZE-1) & MULT_118(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(5)<=signed(MULT_117(5)(MULT_SIZE-1) & MULT_117(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(5)(MULT_SIZE-1) & MULT_118(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(6)<=signed(MULT_117(6)(MULT_SIZE-1) & MULT_117(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(6)(MULT_SIZE-1) & MULT_118(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(7)<=signed(MULT_117(7)(MULT_SIZE-1) & MULT_117(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(7)(MULT_SIZE-1) & MULT_118(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(8)<=signed(MULT_117(8)(MULT_SIZE-1) & MULT_117(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(8)(MULT_SIZE-1) & MULT_118(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(9)<=signed(MULT_117(9)(MULT_SIZE-1) & MULT_117(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(9)(MULT_SIZE-1) & MULT_118(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(10)<=signed(MULT_117(10)(MULT_SIZE-1) & MULT_117(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(10)(MULT_SIZE-1) & MULT_118(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(11)<=signed(MULT_117(11)(MULT_SIZE-1) & MULT_117(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(11)(MULT_SIZE-1) & MULT_118(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(12)<=signed(MULT_117(12)(MULT_SIZE-1) & MULT_117(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(12)(MULT_SIZE-1) & MULT_118(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(13)<=signed(MULT_117(13)(MULT_SIZE-1) & MULT_117(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(13)(MULT_SIZE-1) & MULT_118(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(14)<=signed(MULT_117(14)(MULT_SIZE-1) & MULT_117(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(14)(MULT_SIZE-1) & MULT_118(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(15)<=signed(MULT_117(15)(MULT_SIZE-1) & MULT_117(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(15)(MULT_SIZE-1) & MULT_118(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(16)<=signed(MULT_117(16)(MULT_SIZE-1) & MULT_117(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(16)(MULT_SIZE-1) & MULT_118(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(17)<=signed(MULT_117(17)(MULT_SIZE-1) & MULT_117(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(17)(MULT_SIZE-1) & MULT_118(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(18)<=signed(MULT_117(18)(MULT_SIZE-1) & MULT_117(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(18)(MULT_SIZE-1) & MULT_118(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(19)<=signed(MULT_117(19)(MULT_SIZE-1) & MULT_117(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(19)(MULT_SIZE-1) & MULT_118(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(20)<=signed(MULT_117(20)(MULT_SIZE-1) & MULT_117(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(20)(MULT_SIZE-1) & MULT_118(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(21)<=signed(MULT_117(21)(MULT_SIZE-1) & MULT_117(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(21)(MULT_SIZE-1) & MULT_118(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(22)<=signed(MULT_117(22)(MULT_SIZE-1) & MULT_117(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(22)(MULT_SIZE-1) & MULT_118(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(23)<=signed(MULT_117(23)(MULT_SIZE-1) & MULT_117(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(23)(MULT_SIZE-1) & MULT_118(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(24)<=signed(MULT_117(24)(MULT_SIZE-1) & MULT_117(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(24)(MULT_SIZE-1) & MULT_118(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(25)<=signed(MULT_117(25)(MULT_SIZE-1) & MULT_117(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(25)(MULT_SIZE-1) & MULT_118(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(26)<=signed(MULT_117(26)(MULT_SIZE-1) & MULT_117(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(26)(MULT_SIZE-1) & MULT_118(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(27)<=signed(MULT_117(27)(MULT_SIZE-1) & MULT_117(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(27)(MULT_SIZE-1) & MULT_118(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(28)<=signed(MULT_117(28)(MULT_SIZE-1) & MULT_117(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(28)(MULT_SIZE-1) & MULT_118(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(29)<=signed(MULT_117(29)(MULT_SIZE-1) & MULT_117(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(29)(MULT_SIZE-1) & MULT_118(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(30)<=signed(MULT_117(30)(MULT_SIZE-1) & MULT_117(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(30)(MULT_SIZE-1) & MULT_118(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(31)<=signed(MULT_117(31)(MULT_SIZE-1) & MULT_117(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(31)(MULT_SIZE-1) & MULT_118(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(32)<=signed(MULT_117(32)(MULT_SIZE-1) & MULT_117(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(32)(MULT_SIZE-1) & MULT_118(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(33)<=signed(MULT_117(33)(MULT_SIZE-1) & MULT_117(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(33)(MULT_SIZE-1) & MULT_118(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(34)<=signed(MULT_117(34)(MULT_SIZE-1) & MULT_117(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(34)(MULT_SIZE-1) & MULT_118(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(35)<=signed(MULT_117(35)(MULT_SIZE-1) & MULT_117(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(35)(MULT_SIZE-1) & MULT_118(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(36)<=signed(MULT_117(36)(MULT_SIZE-1) & MULT_117(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(36)(MULT_SIZE-1) & MULT_118(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(37)<=signed(MULT_117(37)(MULT_SIZE-1) & MULT_117(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(37)(MULT_SIZE-1) & MULT_118(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(38)<=signed(MULT_117(38)(MULT_SIZE-1) & MULT_117(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(38)(MULT_SIZE-1) & MULT_118(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(39)<=signed(MULT_117(39)(MULT_SIZE-1) & MULT_117(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(39)(MULT_SIZE-1) & MULT_118(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(40)<=signed(MULT_117(40)(MULT_SIZE-1) & MULT_117(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(40)(MULT_SIZE-1) & MULT_118(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(41)<=signed(MULT_117(41)(MULT_SIZE-1) & MULT_117(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(41)(MULT_SIZE-1) & MULT_118(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(42)<=signed(MULT_117(42)(MULT_SIZE-1) & MULT_117(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(42)(MULT_SIZE-1) & MULT_118(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(43)<=signed(MULT_117(43)(MULT_SIZE-1) & MULT_117(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(43)(MULT_SIZE-1) & MULT_118(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(44)<=signed(MULT_117(44)(MULT_SIZE-1) & MULT_117(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(44)(MULT_SIZE-1) & MULT_118(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(45)<=signed(MULT_117(45)(MULT_SIZE-1) & MULT_117(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(45)(MULT_SIZE-1) & MULT_118(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(46)<=signed(MULT_117(46)(MULT_SIZE-1) & MULT_117(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(46)(MULT_SIZE-1) & MULT_118(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(47)<=signed(MULT_117(47)(MULT_SIZE-1) & MULT_117(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(47)(MULT_SIZE-1) & MULT_118(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(48)<=signed(MULT_117(48)(MULT_SIZE-1) & MULT_117(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(48)(MULT_SIZE-1) & MULT_118(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(49)<=signed(MULT_117(49)(MULT_SIZE-1) & MULT_117(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(49)(MULT_SIZE-1) & MULT_118(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(50)<=signed(MULT_117(50)(MULT_SIZE-1) & MULT_117(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(50)(MULT_SIZE-1) & MULT_118(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(51)<=signed(MULT_117(51)(MULT_SIZE-1) & MULT_117(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(51)(MULT_SIZE-1) & MULT_118(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(52)<=signed(MULT_117(52)(MULT_SIZE-1) & MULT_117(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(52)(MULT_SIZE-1) & MULT_118(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(53)<=signed(MULT_117(53)(MULT_SIZE-1) & MULT_117(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(53)(MULT_SIZE-1) & MULT_118(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(54)<=signed(MULT_117(54)(MULT_SIZE-1) & MULT_117(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(54)(MULT_SIZE-1) & MULT_118(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(55)<=signed(MULT_117(55)(MULT_SIZE-1) & MULT_117(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(55)(MULT_SIZE-1) & MULT_118(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(56)<=signed(MULT_117(56)(MULT_SIZE-1) & MULT_117(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(56)(MULT_SIZE-1) & MULT_118(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(57)<=signed(MULT_117(57)(MULT_SIZE-1) & MULT_117(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(57)(MULT_SIZE-1) & MULT_118(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(58)<=signed(MULT_117(58)(MULT_SIZE-1) & MULT_117(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(58)(MULT_SIZE-1) & MULT_118(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(59)<=signed(MULT_117(59)(MULT_SIZE-1) & MULT_117(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(59)(MULT_SIZE-1) & MULT_118(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(60)<=signed(MULT_117(60)(MULT_SIZE-1) & MULT_117(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(60)(MULT_SIZE-1) & MULT_118(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(61)<=signed(MULT_117(61)(MULT_SIZE-1) & MULT_117(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(61)(MULT_SIZE-1) & MULT_118(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(62)<=signed(MULT_117(62)(MULT_SIZE-1) & MULT_117(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(62)(MULT_SIZE-1) & MULT_118(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(63)<=signed(MULT_117(63)(MULT_SIZE-1) & MULT_117(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(63)(MULT_SIZE-1) & MULT_118(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(64)<=signed(MULT_117(64)(MULT_SIZE-1) & MULT_117(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(64)(MULT_SIZE-1) & MULT_118(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(65)<=signed(MULT_117(65)(MULT_SIZE-1) & MULT_117(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(65)(MULT_SIZE-1) & MULT_118(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(66)<=signed(MULT_117(66)(MULT_SIZE-1) & MULT_117(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(66)(MULT_SIZE-1) & MULT_118(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(67)<=signed(MULT_117(67)(MULT_SIZE-1) & MULT_117(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(67)(MULT_SIZE-1) & MULT_118(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(68)<=signed(MULT_117(68)(MULT_SIZE-1) & MULT_117(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(68)(MULT_SIZE-1) & MULT_118(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(69)<=signed(MULT_117(69)(MULT_SIZE-1) & MULT_117(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(69)(MULT_SIZE-1) & MULT_118(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(70)<=signed(MULT_117(70)(MULT_SIZE-1) & MULT_117(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(70)(MULT_SIZE-1) & MULT_118(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(71)<=signed(MULT_117(71)(MULT_SIZE-1) & MULT_117(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(71)(MULT_SIZE-1) & MULT_118(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(72)<=signed(MULT_117(72)(MULT_SIZE-1) & MULT_117(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(72)(MULT_SIZE-1) & MULT_118(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(73)<=signed(MULT_117(73)(MULT_SIZE-1) & MULT_117(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(73)(MULT_SIZE-1) & MULT_118(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(74)<=signed(MULT_117(74)(MULT_SIZE-1) & MULT_117(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(74)(MULT_SIZE-1) & MULT_118(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(75)<=signed(MULT_117(75)(MULT_SIZE-1) & MULT_117(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(75)(MULT_SIZE-1) & MULT_118(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(76)<=signed(MULT_117(76)(MULT_SIZE-1) & MULT_117(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(76)(MULT_SIZE-1) & MULT_118(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(77)<=signed(MULT_117(77)(MULT_SIZE-1) & MULT_117(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(77)(MULT_SIZE-1) & MULT_118(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(78)<=signed(MULT_117(78)(MULT_SIZE-1) & MULT_117(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(78)(MULT_SIZE-1) & MULT_118(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(79)<=signed(MULT_117(79)(MULT_SIZE-1) & MULT_117(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(79)(MULT_SIZE-1) & MULT_118(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(80)<=signed(MULT_117(80)(MULT_SIZE-1) & MULT_117(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(80)(MULT_SIZE-1) & MULT_118(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(81)<=signed(MULT_117(81)(MULT_SIZE-1) & MULT_117(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(81)(MULT_SIZE-1) & MULT_118(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(82)<=signed(MULT_117(82)(MULT_SIZE-1) & MULT_117(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(82)(MULT_SIZE-1) & MULT_118(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_59(83)<=signed(MULT_117(83)(MULT_SIZE-1) & MULT_117(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_118(83)(MULT_SIZE-1) & MULT_118(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));

			MULTS_1_60(0)<=signed(MULT_119(0)(MULT_SIZE-1) & MULT_119(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(0)(MULT_SIZE-1) & MULT_120(0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(1)<=signed(MULT_119(1)(MULT_SIZE-1) & MULT_119(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(1)(MULT_SIZE-1) & MULT_120(1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(2)<=signed(MULT_119(2)(MULT_SIZE-1) & MULT_119(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(2)(MULT_SIZE-1) & MULT_120(2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(3)<=signed(MULT_119(3)(MULT_SIZE-1) & MULT_119(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(3)(MULT_SIZE-1) & MULT_120(3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(4)<=signed(MULT_119(4)(MULT_SIZE-1) & MULT_119(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(4)(MULT_SIZE-1) & MULT_120(4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(5)<=signed(MULT_119(5)(MULT_SIZE-1) & MULT_119(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(5)(MULT_SIZE-1) & MULT_120(5)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(6)<=signed(MULT_119(6)(MULT_SIZE-1) & MULT_119(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(6)(MULT_SIZE-1) & MULT_120(6)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(7)<=signed(MULT_119(7)(MULT_SIZE-1) & MULT_119(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(7)(MULT_SIZE-1) & MULT_120(7)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(8)<=signed(MULT_119(8)(MULT_SIZE-1) & MULT_119(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(8)(MULT_SIZE-1) & MULT_120(8)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(9)<=signed(MULT_119(9)(MULT_SIZE-1) & MULT_119(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(9)(MULT_SIZE-1) & MULT_120(9)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(10)<=signed(MULT_119(10)(MULT_SIZE-1) & MULT_119(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(10)(MULT_SIZE-1) & MULT_120(10)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(11)<=signed(MULT_119(11)(MULT_SIZE-1) & MULT_119(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(11)(MULT_SIZE-1) & MULT_120(11)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(12)<=signed(MULT_119(12)(MULT_SIZE-1) & MULT_119(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(12)(MULT_SIZE-1) & MULT_120(12)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(13)<=signed(MULT_119(13)(MULT_SIZE-1) & MULT_119(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(13)(MULT_SIZE-1) & MULT_120(13)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(14)<=signed(MULT_119(14)(MULT_SIZE-1) & MULT_119(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(14)(MULT_SIZE-1) & MULT_120(14)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(15)<=signed(MULT_119(15)(MULT_SIZE-1) & MULT_119(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(15)(MULT_SIZE-1) & MULT_120(15)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(16)<=signed(MULT_119(16)(MULT_SIZE-1) & MULT_119(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(16)(MULT_SIZE-1) & MULT_120(16)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(17)<=signed(MULT_119(17)(MULT_SIZE-1) & MULT_119(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(17)(MULT_SIZE-1) & MULT_120(17)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(18)<=signed(MULT_119(18)(MULT_SIZE-1) & MULT_119(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(18)(MULT_SIZE-1) & MULT_120(18)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(19)<=signed(MULT_119(19)(MULT_SIZE-1) & MULT_119(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(19)(MULT_SIZE-1) & MULT_120(19)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(20)<=signed(MULT_119(20)(MULT_SIZE-1) & MULT_119(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(20)(MULT_SIZE-1) & MULT_120(20)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(21)<=signed(MULT_119(21)(MULT_SIZE-1) & MULT_119(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(21)(MULT_SIZE-1) & MULT_120(21)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(22)<=signed(MULT_119(22)(MULT_SIZE-1) & MULT_119(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(22)(MULT_SIZE-1) & MULT_120(22)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(23)<=signed(MULT_119(23)(MULT_SIZE-1) & MULT_119(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(23)(MULT_SIZE-1) & MULT_120(23)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(24)<=signed(MULT_119(24)(MULT_SIZE-1) & MULT_119(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(24)(MULT_SIZE-1) & MULT_120(24)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(25)<=signed(MULT_119(25)(MULT_SIZE-1) & MULT_119(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(25)(MULT_SIZE-1) & MULT_120(25)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(26)<=signed(MULT_119(26)(MULT_SIZE-1) & MULT_119(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(26)(MULT_SIZE-1) & MULT_120(26)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(27)<=signed(MULT_119(27)(MULT_SIZE-1) & MULT_119(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(27)(MULT_SIZE-1) & MULT_120(27)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(28)<=signed(MULT_119(28)(MULT_SIZE-1) & MULT_119(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(28)(MULT_SIZE-1) & MULT_120(28)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(29)<=signed(MULT_119(29)(MULT_SIZE-1) & MULT_119(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(29)(MULT_SIZE-1) & MULT_120(29)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(30)<=signed(MULT_119(30)(MULT_SIZE-1) & MULT_119(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(30)(MULT_SIZE-1) & MULT_120(30)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(31)<=signed(MULT_119(31)(MULT_SIZE-1) & MULT_119(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(31)(MULT_SIZE-1) & MULT_120(31)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(32)<=signed(MULT_119(32)(MULT_SIZE-1) & MULT_119(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(32)(MULT_SIZE-1) & MULT_120(32)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(33)<=signed(MULT_119(33)(MULT_SIZE-1) & MULT_119(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(33)(MULT_SIZE-1) & MULT_120(33)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(34)<=signed(MULT_119(34)(MULT_SIZE-1) & MULT_119(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(34)(MULT_SIZE-1) & MULT_120(34)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(35)<=signed(MULT_119(35)(MULT_SIZE-1) & MULT_119(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(35)(MULT_SIZE-1) & MULT_120(35)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(36)<=signed(MULT_119(36)(MULT_SIZE-1) & MULT_119(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(36)(MULT_SIZE-1) & MULT_120(36)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(37)<=signed(MULT_119(37)(MULT_SIZE-1) & MULT_119(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(37)(MULT_SIZE-1) & MULT_120(37)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(38)<=signed(MULT_119(38)(MULT_SIZE-1) & MULT_119(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(38)(MULT_SIZE-1) & MULT_120(38)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(39)<=signed(MULT_119(39)(MULT_SIZE-1) & MULT_119(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(39)(MULT_SIZE-1) & MULT_120(39)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(40)<=signed(MULT_119(40)(MULT_SIZE-1) & MULT_119(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(40)(MULT_SIZE-1) & MULT_120(40)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(41)<=signed(MULT_119(41)(MULT_SIZE-1) & MULT_119(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(41)(MULT_SIZE-1) & MULT_120(41)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(42)<=signed(MULT_119(42)(MULT_SIZE-1) & MULT_119(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(42)(MULT_SIZE-1) & MULT_120(42)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(43)<=signed(MULT_119(43)(MULT_SIZE-1) & MULT_119(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(43)(MULT_SIZE-1) & MULT_120(43)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(44)<=signed(MULT_119(44)(MULT_SIZE-1) & MULT_119(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(44)(MULT_SIZE-1) & MULT_120(44)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(45)<=signed(MULT_119(45)(MULT_SIZE-1) & MULT_119(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(45)(MULT_SIZE-1) & MULT_120(45)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(46)<=signed(MULT_119(46)(MULT_SIZE-1) & MULT_119(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(46)(MULT_SIZE-1) & MULT_120(46)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(47)<=signed(MULT_119(47)(MULT_SIZE-1) & MULT_119(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(47)(MULT_SIZE-1) & MULT_120(47)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(48)<=signed(MULT_119(48)(MULT_SIZE-1) & MULT_119(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(48)(MULT_SIZE-1) & MULT_120(48)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(49)<=signed(MULT_119(49)(MULT_SIZE-1) & MULT_119(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(49)(MULT_SIZE-1) & MULT_120(49)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(50)<=signed(MULT_119(50)(MULT_SIZE-1) & MULT_119(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(50)(MULT_SIZE-1) & MULT_120(50)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(51)<=signed(MULT_119(51)(MULT_SIZE-1) & MULT_119(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(51)(MULT_SIZE-1) & MULT_120(51)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(52)<=signed(MULT_119(52)(MULT_SIZE-1) & MULT_119(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(52)(MULT_SIZE-1) & MULT_120(52)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(53)<=signed(MULT_119(53)(MULT_SIZE-1) & MULT_119(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(53)(MULT_SIZE-1) & MULT_120(53)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(54)<=signed(MULT_119(54)(MULT_SIZE-1) & MULT_119(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(54)(MULT_SIZE-1) & MULT_120(54)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(55)<=signed(MULT_119(55)(MULT_SIZE-1) & MULT_119(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(55)(MULT_SIZE-1) & MULT_120(55)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(56)<=signed(MULT_119(56)(MULT_SIZE-1) & MULT_119(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(56)(MULT_SIZE-1) & MULT_120(56)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(57)<=signed(MULT_119(57)(MULT_SIZE-1) & MULT_119(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(57)(MULT_SIZE-1) & MULT_120(57)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(58)<=signed(MULT_119(58)(MULT_SIZE-1) & MULT_119(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(58)(MULT_SIZE-1) & MULT_120(58)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(59)<=signed(MULT_119(59)(MULT_SIZE-1) & MULT_119(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(59)(MULT_SIZE-1) & MULT_120(59)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(60)<=signed(MULT_119(60)(MULT_SIZE-1) & MULT_119(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(60)(MULT_SIZE-1) & MULT_120(60)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(61)<=signed(MULT_119(61)(MULT_SIZE-1) & MULT_119(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(61)(MULT_SIZE-1) & MULT_120(61)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(62)<=signed(MULT_119(62)(MULT_SIZE-1) & MULT_119(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(62)(MULT_SIZE-1) & MULT_120(62)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(63)<=signed(MULT_119(63)(MULT_SIZE-1) & MULT_119(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(63)(MULT_SIZE-1) & MULT_120(63)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(64)<=signed(MULT_119(64)(MULT_SIZE-1) & MULT_119(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(64)(MULT_SIZE-1) & MULT_120(64)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(65)<=signed(MULT_119(65)(MULT_SIZE-1) & MULT_119(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(65)(MULT_SIZE-1) & MULT_120(65)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(66)<=signed(MULT_119(66)(MULT_SIZE-1) & MULT_119(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(66)(MULT_SIZE-1) & MULT_120(66)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(67)<=signed(MULT_119(67)(MULT_SIZE-1) & MULT_119(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(67)(MULT_SIZE-1) & MULT_120(67)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(68)<=signed(MULT_119(68)(MULT_SIZE-1) & MULT_119(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(68)(MULT_SIZE-1) & MULT_120(68)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(69)<=signed(MULT_119(69)(MULT_SIZE-1) & MULT_119(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(69)(MULT_SIZE-1) & MULT_120(69)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(70)<=signed(MULT_119(70)(MULT_SIZE-1) & MULT_119(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(70)(MULT_SIZE-1) & MULT_120(70)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(71)<=signed(MULT_119(71)(MULT_SIZE-1) & MULT_119(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(71)(MULT_SIZE-1) & MULT_120(71)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(72)<=signed(MULT_119(72)(MULT_SIZE-1) & MULT_119(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(72)(MULT_SIZE-1) & MULT_120(72)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(73)<=signed(MULT_119(73)(MULT_SIZE-1) & MULT_119(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(73)(MULT_SIZE-1) & MULT_120(73)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(74)<=signed(MULT_119(74)(MULT_SIZE-1) & MULT_119(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(74)(MULT_SIZE-1) & MULT_120(74)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(75)<=signed(MULT_119(75)(MULT_SIZE-1) & MULT_119(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(75)(MULT_SIZE-1) & MULT_120(75)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(76)<=signed(MULT_119(76)(MULT_SIZE-1) & MULT_119(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(76)(MULT_SIZE-1) & MULT_120(76)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(77)<=signed(MULT_119(77)(MULT_SIZE-1) & MULT_119(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(77)(MULT_SIZE-1) & MULT_120(77)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(78)<=signed(MULT_119(78)(MULT_SIZE-1) & MULT_119(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(78)(MULT_SIZE-1) & MULT_120(78)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(79)<=signed(MULT_119(79)(MULT_SIZE-1) & MULT_119(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(79)(MULT_SIZE-1) & MULT_120(79)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(80)<=signed(MULT_119(80)(MULT_SIZE-1) & MULT_119(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(80)(MULT_SIZE-1) & MULT_120(80)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(81)<=signed(MULT_119(81)(MULT_SIZE-1) & MULT_119(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(81)(MULT_SIZE-1) & MULT_120(81)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(82)<=signed(MULT_119(82)(MULT_SIZE-1) & MULT_119(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(82)(MULT_SIZE-1) & MULT_120(82)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_60(83)<=signed(MULT_119(83)(MULT_SIZE-1) & MULT_119(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2))+signed(MULT_120(83)(MULT_SIZE-1) & MULT_120(83)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));



                     EN_SUM_MULT_2<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_2 = '1' then
			------------------------------------STAGE-2--------------------------------------
			MULTS_2_1(0)<=signed(MULTS_1_1(0)(PERCISION) & MULTS_1_1(0)(PERCISION downto 1))+signed(MULTS_1_2(0)(PERCISION) & MULTS_1_2(0)(PERCISION downto 1));
			MULTS_2_1(1)<=signed(MULTS_1_1(1)(PERCISION) & MULTS_1_1(1)(PERCISION downto 1))+signed(MULTS_1_2(1)(PERCISION) & MULTS_1_2(1)(PERCISION downto 1));
			MULTS_2_1(2)<=signed(MULTS_1_1(2)(PERCISION) & MULTS_1_1(2)(PERCISION downto 1))+signed(MULTS_1_2(2)(PERCISION) & MULTS_1_2(2)(PERCISION downto 1));
			MULTS_2_1(3)<=signed(MULTS_1_1(3)(PERCISION) & MULTS_1_1(3)(PERCISION downto 1))+signed(MULTS_1_2(3)(PERCISION) & MULTS_1_2(3)(PERCISION downto 1));
			MULTS_2_1(4)<=signed(MULTS_1_1(4)(PERCISION) & MULTS_1_1(4)(PERCISION downto 1))+signed(MULTS_1_2(4)(PERCISION) & MULTS_1_2(4)(PERCISION downto 1));
			MULTS_2_1(5)<=signed(MULTS_1_1(5)(PERCISION) & MULTS_1_1(5)(PERCISION downto 1))+signed(MULTS_1_2(5)(PERCISION) & MULTS_1_2(5)(PERCISION downto 1));
			MULTS_2_1(6)<=signed(MULTS_1_1(6)(PERCISION) & MULTS_1_1(6)(PERCISION downto 1))+signed(MULTS_1_2(6)(PERCISION) & MULTS_1_2(6)(PERCISION downto 1));
			MULTS_2_1(7)<=signed(MULTS_1_1(7)(PERCISION) & MULTS_1_1(7)(PERCISION downto 1))+signed(MULTS_1_2(7)(PERCISION) & MULTS_1_2(7)(PERCISION downto 1));
			MULTS_2_1(8)<=signed(MULTS_1_1(8)(PERCISION) & MULTS_1_1(8)(PERCISION downto 1))+signed(MULTS_1_2(8)(PERCISION) & MULTS_1_2(8)(PERCISION downto 1));
			MULTS_2_1(9)<=signed(MULTS_1_1(9)(PERCISION) & MULTS_1_1(9)(PERCISION downto 1))+signed(MULTS_1_2(9)(PERCISION) & MULTS_1_2(9)(PERCISION downto 1));
			MULTS_2_1(10)<=signed(MULTS_1_1(10)(PERCISION) & MULTS_1_1(10)(PERCISION downto 1))+signed(MULTS_1_2(10)(PERCISION) & MULTS_1_2(10)(PERCISION downto 1));
			MULTS_2_1(11)<=signed(MULTS_1_1(11)(PERCISION) & MULTS_1_1(11)(PERCISION downto 1))+signed(MULTS_1_2(11)(PERCISION) & MULTS_1_2(11)(PERCISION downto 1));
			MULTS_2_1(12)<=signed(MULTS_1_1(12)(PERCISION) & MULTS_1_1(12)(PERCISION downto 1))+signed(MULTS_1_2(12)(PERCISION) & MULTS_1_2(12)(PERCISION downto 1));
			MULTS_2_1(13)<=signed(MULTS_1_1(13)(PERCISION) & MULTS_1_1(13)(PERCISION downto 1))+signed(MULTS_1_2(13)(PERCISION) & MULTS_1_2(13)(PERCISION downto 1));
			MULTS_2_1(14)<=signed(MULTS_1_1(14)(PERCISION) & MULTS_1_1(14)(PERCISION downto 1))+signed(MULTS_1_2(14)(PERCISION) & MULTS_1_2(14)(PERCISION downto 1));
			MULTS_2_1(15)<=signed(MULTS_1_1(15)(PERCISION) & MULTS_1_1(15)(PERCISION downto 1))+signed(MULTS_1_2(15)(PERCISION) & MULTS_1_2(15)(PERCISION downto 1));
			MULTS_2_1(16)<=signed(MULTS_1_1(16)(PERCISION) & MULTS_1_1(16)(PERCISION downto 1))+signed(MULTS_1_2(16)(PERCISION) & MULTS_1_2(16)(PERCISION downto 1));
			MULTS_2_1(17)<=signed(MULTS_1_1(17)(PERCISION) & MULTS_1_1(17)(PERCISION downto 1))+signed(MULTS_1_2(17)(PERCISION) & MULTS_1_2(17)(PERCISION downto 1));
			MULTS_2_1(18)<=signed(MULTS_1_1(18)(PERCISION) & MULTS_1_1(18)(PERCISION downto 1))+signed(MULTS_1_2(18)(PERCISION) & MULTS_1_2(18)(PERCISION downto 1));
			MULTS_2_1(19)<=signed(MULTS_1_1(19)(PERCISION) & MULTS_1_1(19)(PERCISION downto 1))+signed(MULTS_1_2(19)(PERCISION) & MULTS_1_2(19)(PERCISION downto 1));
			MULTS_2_1(20)<=signed(MULTS_1_1(20)(PERCISION) & MULTS_1_1(20)(PERCISION downto 1))+signed(MULTS_1_2(20)(PERCISION) & MULTS_1_2(20)(PERCISION downto 1));
			MULTS_2_1(21)<=signed(MULTS_1_1(21)(PERCISION) & MULTS_1_1(21)(PERCISION downto 1))+signed(MULTS_1_2(21)(PERCISION) & MULTS_1_2(21)(PERCISION downto 1));
			MULTS_2_1(22)<=signed(MULTS_1_1(22)(PERCISION) & MULTS_1_1(22)(PERCISION downto 1))+signed(MULTS_1_2(22)(PERCISION) & MULTS_1_2(22)(PERCISION downto 1));
			MULTS_2_1(23)<=signed(MULTS_1_1(23)(PERCISION) & MULTS_1_1(23)(PERCISION downto 1))+signed(MULTS_1_2(23)(PERCISION) & MULTS_1_2(23)(PERCISION downto 1));
			MULTS_2_1(24)<=signed(MULTS_1_1(24)(PERCISION) & MULTS_1_1(24)(PERCISION downto 1))+signed(MULTS_1_2(24)(PERCISION) & MULTS_1_2(24)(PERCISION downto 1));
			MULTS_2_1(25)<=signed(MULTS_1_1(25)(PERCISION) & MULTS_1_1(25)(PERCISION downto 1))+signed(MULTS_1_2(25)(PERCISION) & MULTS_1_2(25)(PERCISION downto 1));
			MULTS_2_1(26)<=signed(MULTS_1_1(26)(PERCISION) & MULTS_1_1(26)(PERCISION downto 1))+signed(MULTS_1_2(26)(PERCISION) & MULTS_1_2(26)(PERCISION downto 1));
			MULTS_2_1(27)<=signed(MULTS_1_1(27)(PERCISION) & MULTS_1_1(27)(PERCISION downto 1))+signed(MULTS_1_2(27)(PERCISION) & MULTS_1_2(27)(PERCISION downto 1));
			MULTS_2_1(28)<=signed(MULTS_1_1(28)(PERCISION) & MULTS_1_1(28)(PERCISION downto 1))+signed(MULTS_1_2(28)(PERCISION) & MULTS_1_2(28)(PERCISION downto 1));
			MULTS_2_1(29)<=signed(MULTS_1_1(29)(PERCISION) & MULTS_1_1(29)(PERCISION downto 1))+signed(MULTS_1_2(29)(PERCISION) & MULTS_1_2(29)(PERCISION downto 1));
			MULTS_2_1(30)<=signed(MULTS_1_1(30)(PERCISION) & MULTS_1_1(30)(PERCISION downto 1))+signed(MULTS_1_2(30)(PERCISION) & MULTS_1_2(30)(PERCISION downto 1));
			MULTS_2_1(31)<=signed(MULTS_1_1(31)(PERCISION) & MULTS_1_1(31)(PERCISION downto 1))+signed(MULTS_1_2(31)(PERCISION) & MULTS_1_2(31)(PERCISION downto 1));
			MULTS_2_1(32)<=signed(MULTS_1_1(32)(PERCISION) & MULTS_1_1(32)(PERCISION downto 1))+signed(MULTS_1_2(32)(PERCISION) & MULTS_1_2(32)(PERCISION downto 1));
			MULTS_2_1(33)<=signed(MULTS_1_1(33)(PERCISION) & MULTS_1_1(33)(PERCISION downto 1))+signed(MULTS_1_2(33)(PERCISION) & MULTS_1_2(33)(PERCISION downto 1));
			MULTS_2_1(34)<=signed(MULTS_1_1(34)(PERCISION) & MULTS_1_1(34)(PERCISION downto 1))+signed(MULTS_1_2(34)(PERCISION) & MULTS_1_2(34)(PERCISION downto 1));
			MULTS_2_1(35)<=signed(MULTS_1_1(35)(PERCISION) & MULTS_1_1(35)(PERCISION downto 1))+signed(MULTS_1_2(35)(PERCISION) & MULTS_1_2(35)(PERCISION downto 1));
			MULTS_2_1(36)<=signed(MULTS_1_1(36)(PERCISION) & MULTS_1_1(36)(PERCISION downto 1))+signed(MULTS_1_2(36)(PERCISION) & MULTS_1_2(36)(PERCISION downto 1));
			MULTS_2_1(37)<=signed(MULTS_1_1(37)(PERCISION) & MULTS_1_1(37)(PERCISION downto 1))+signed(MULTS_1_2(37)(PERCISION) & MULTS_1_2(37)(PERCISION downto 1));
			MULTS_2_1(38)<=signed(MULTS_1_1(38)(PERCISION) & MULTS_1_1(38)(PERCISION downto 1))+signed(MULTS_1_2(38)(PERCISION) & MULTS_1_2(38)(PERCISION downto 1));
			MULTS_2_1(39)<=signed(MULTS_1_1(39)(PERCISION) & MULTS_1_1(39)(PERCISION downto 1))+signed(MULTS_1_2(39)(PERCISION) & MULTS_1_2(39)(PERCISION downto 1));
			MULTS_2_1(40)<=signed(MULTS_1_1(40)(PERCISION) & MULTS_1_1(40)(PERCISION downto 1))+signed(MULTS_1_2(40)(PERCISION) & MULTS_1_2(40)(PERCISION downto 1));
			MULTS_2_1(41)<=signed(MULTS_1_1(41)(PERCISION) & MULTS_1_1(41)(PERCISION downto 1))+signed(MULTS_1_2(41)(PERCISION) & MULTS_1_2(41)(PERCISION downto 1));
			MULTS_2_1(42)<=signed(MULTS_1_1(42)(PERCISION) & MULTS_1_1(42)(PERCISION downto 1))+signed(MULTS_1_2(42)(PERCISION) & MULTS_1_2(42)(PERCISION downto 1));
			MULTS_2_1(43)<=signed(MULTS_1_1(43)(PERCISION) & MULTS_1_1(43)(PERCISION downto 1))+signed(MULTS_1_2(43)(PERCISION) & MULTS_1_2(43)(PERCISION downto 1));
			MULTS_2_1(44)<=signed(MULTS_1_1(44)(PERCISION) & MULTS_1_1(44)(PERCISION downto 1))+signed(MULTS_1_2(44)(PERCISION) & MULTS_1_2(44)(PERCISION downto 1));
			MULTS_2_1(45)<=signed(MULTS_1_1(45)(PERCISION) & MULTS_1_1(45)(PERCISION downto 1))+signed(MULTS_1_2(45)(PERCISION) & MULTS_1_2(45)(PERCISION downto 1));
			MULTS_2_1(46)<=signed(MULTS_1_1(46)(PERCISION) & MULTS_1_1(46)(PERCISION downto 1))+signed(MULTS_1_2(46)(PERCISION) & MULTS_1_2(46)(PERCISION downto 1));
			MULTS_2_1(47)<=signed(MULTS_1_1(47)(PERCISION) & MULTS_1_1(47)(PERCISION downto 1))+signed(MULTS_1_2(47)(PERCISION) & MULTS_1_2(47)(PERCISION downto 1));
			MULTS_2_1(48)<=signed(MULTS_1_1(48)(PERCISION) & MULTS_1_1(48)(PERCISION downto 1))+signed(MULTS_1_2(48)(PERCISION) & MULTS_1_2(48)(PERCISION downto 1));
			MULTS_2_1(49)<=signed(MULTS_1_1(49)(PERCISION) & MULTS_1_1(49)(PERCISION downto 1))+signed(MULTS_1_2(49)(PERCISION) & MULTS_1_2(49)(PERCISION downto 1));
			MULTS_2_1(50)<=signed(MULTS_1_1(50)(PERCISION) & MULTS_1_1(50)(PERCISION downto 1))+signed(MULTS_1_2(50)(PERCISION) & MULTS_1_2(50)(PERCISION downto 1));
			MULTS_2_1(51)<=signed(MULTS_1_1(51)(PERCISION) & MULTS_1_1(51)(PERCISION downto 1))+signed(MULTS_1_2(51)(PERCISION) & MULTS_1_2(51)(PERCISION downto 1));
			MULTS_2_1(52)<=signed(MULTS_1_1(52)(PERCISION) & MULTS_1_1(52)(PERCISION downto 1))+signed(MULTS_1_2(52)(PERCISION) & MULTS_1_2(52)(PERCISION downto 1));
			MULTS_2_1(53)<=signed(MULTS_1_1(53)(PERCISION) & MULTS_1_1(53)(PERCISION downto 1))+signed(MULTS_1_2(53)(PERCISION) & MULTS_1_2(53)(PERCISION downto 1));
			MULTS_2_1(54)<=signed(MULTS_1_1(54)(PERCISION) & MULTS_1_1(54)(PERCISION downto 1))+signed(MULTS_1_2(54)(PERCISION) & MULTS_1_2(54)(PERCISION downto 1));
			MULTS_2_1(55)<=signed(MULTS_1_1(55)(PERCISION) & MULTS_1_1(55)(PERCISION downto 1))+signed(MULTS_1_2(55)(PERCISION) & MULTS_1_2(55)(PERCISION downto 1));
			MULTS_2_1(56)<=signed(MULTS_1_1(56)(PERCISION) & MULTS_1_1(56)(PERCISION downto 1))+signed(MULTS_1_2(56)(PERCISION) & MULTS_1_2(56)(PERCISION downto 1));
			MULTS_2_1(57)<=signed(MULTS_1_1(57)(PERCISION) & MULTS_1_1(57)(PERCISION downto 1))+signed(MULTS_1_2(57)(PERCISION) & MULTS_1_2(57)(PERCISION downto 1));
			MULTS_2_1(58)<=signed(MULTS_1_1(58)(PERCISION) & MULTS_1_1(58)(PERCISION downto 1))+signed(MULTS_1_2(58)(PERCISION) & MULTS_1_2(58)(PERCISION downto 1));
			MULTS_2_1(59)<=signed(MULTS_1_1(59)(PERCISION) & MULTS_1_1(59)(PERCISION downto 1))+signed(MULTS_1_2(59)(PERCISION) & MULTS_1_2(59)(PERCISION downto 1));
			MULTS_2_1(60)<=signed(MULTS_1_1(60)(PERCISION) & MULTS_1_1(60)(PERCISION downto 1))+signed(MULTS_1_2(60)(PERCISION) & MULTS_1_2(60)(PERCISION downto 1));
			MULTS_2_1(61)<=signed(MULTS_1_1(61)(PERCISION) & MULTS_1_1(61)(PERCISION downto 1))+signed(MULTS_1_2(61)(PERCISION) & MULTS_1_2(61)(PERCISION downto 1));
			MULTS_2_1(62)<=signed(MULTS_1_1(62)(PERCISION) & MULTS_1_1(62)(PERCISION downto 1))+signed(MULTS_1_2(62)(PERCISION) & MULTS_1_2(62)(PERCISION downto 1));
			MULTS_2_1(63)<=signed(MULTS_1_1(63)(PERCISION) & MULTS_1_1(63)(PERCISION downto 1))+signed(MULTS_1_2(63)(PERCISION) & MULTS_1_2(63)(PERCISION downto 1));
			MULTS_2_1(64)<=signed(MULTS_1_1(64)(PERCISION) & MULTS_1_1(64)(PERCISION downto 1))+signed(MULTS_1_2(64)(PERCISION) & MULTS_1_2(64)(PERCISION downto 1));
			MULTS_2_1(65)<=signed(MULTS_1_1(65)(PERCISION) & MULTS_1_1(65)(PERCISION downto 1))+signed(MULTS_1_2(65)(PERCISION) & MULTS_1_2(65)(PERCISION downto 1));
			MULTS_2_1(66)<=signed(MULTS_1_1(66)(PERCISION) & MULTS_1_1(66)(PERCISION downto 1))+signed(MULTS_1_2(66)(PERCISION) & MULTS_1_2(66)(PERCISION downto 1));
			MULTS_2_1(67)<=signed(MULTS_1_1(67)(PERCISION) & MULTS_1_1(67)(PERCISION downto 1))+signed(MULTS_1_2(67)(PERCISION) & MULTS_1_2(67)(PERCISION downto 1));
			MULTS_2_1(68)<=signed(MULTS_1_1(68)(PERCISION) & MULTS_1_1(68)(PERCISION downto 1))+signed(MULTS_1_2(68)(PERCISION) & MULTS_1_2(68)(PERCISION downto 1));
			MULTS_2_1(69)<=signed(MULTS_1_1(69)(PERCISION) & MULTS_1_1(69)(PERCISION downto 1))+signed(MULTS_1_2(69)(PERCISION) & MULTS_1_2(69)(PERCISION downto 1));
			MULTS_2_1(70)<=signed(MULTS_1_1(70)(PERCISION) & MULTS_1_1(70)(PERCISION downto 1))+signed(MULTS_1_2(70)(PERCISION) & MULTS_1_2(70)(PERCISION downto 1));
			MULTS_2_1(71)<=signed(MULTS_1_1(71)(PERCISION) & MULTS_1_1(71)(PERCISION downto 1))+signed(MULTS_1_2(71)(PERCISION) & MULTS_1_2(71)(PERCISION downto 1));
			MULTS_2_1(72)<=signed(MULTS_1_1(72)(PERCISION) & MULTS_1_1(72)(PERCISION downto 1))+signed(MULTS_1_2(72)(PERCISION) & MULTS_1_2(72)(PERCISION downto 1));
			MULTS_2_1(73)<=signed(MULTS_1_1(73)(PERCISION) & MULTS_1_1(73)(PERCISION downto 1))+signed(MULTS_1_2(73)(PERCISION) & MULTS_1_2(73)(PERCISION downto 1));
			MULTS_2_1(74)<=signed(MULTS_1_1(74)(PERCISION) & MULTS_1_1(74)(PERCISION downto 1))+signed(MULTS_1_2(74)(PERCISION) & MULTS_1_2(74)(PERCISION downto 1));
			MULTS_2_1(75)<=signed(MULTS_1_1(75)(PERCISION) & MULTS_1_1(75)(PERCISION downto 1))+signed(MULTS_1_2(75)(PERCISION) & MULTS_1_2(75)(PERCISION downto 1));
			MULTS_2_1(76)<=signed(MULTS_1_1(76)(PERCISION) & MULTS_1_1(76)(PERCISION downto 1))+signed(MULTS_1_2(76)(PERCISION) & MULTS_1_2(76)(PERCISION downto 1));
			MULTS_2_1(77)<=signed(MULTS_1_1(77)(PERCISION) & MULTS_1_1(77)(PERCISION downto 1))+signed(MULTS_1_2(77)(PERCISION) & MULTS_1_2(77)(PERCISION downto 1));
			MULTS_2_1(78)<=signed(MULTS_1_1(78)(PERCISION) & MULTS_1_1(78)(PERCISION downto 1))+signed(MULTS_1_2(78)(PERCISION) & MULTS_1_2(78)(PERCISION downto 1));
			MULTS_2_1(79)<=signed(MULTS_1_1(79)(PERCISION) & MULTS_1_1(79)(PERCISION downto 1))+signed(MULTS_1_2(79)(PERCISION) & MULTS_1_2(79)(PERCISION downto 1));
			MULTS_2_1(80)<=signed(MULTS_1_1(80)(PERCISION) & MULTS_1_1(80)(PERCISION downto 1))+signed(MULTS_1_2(80)(PERCISION) & MULTS_1_2(80)(PERCISION downto 1));
			MULTS_2_1(81)<=signed(MULTS_1_1(81)(PERCISION) & MULTS_1_1(81)(PERCISION downto 1))+signed(MULTS_1_2(81)(PERCISION) & MULTS_1_2(81)(PERCISION downto 1));
			MULTS_2_1(82)<=signed(MULTS_1_1(82)(PERCISION) & MULTS_1_1(82)(PERCISION downto 1))+signed(MULTS_1_2(82)(PERCISION) & MULTS_1_2(82)(PERCISION downto 1));
			MULTS_2_1(83)<=signed(MULTS_1_1(83)(PERCISION) & MULTS_1_1(83)(PERCISION downto 1))+signed(MULTS_1_2(83)(PERCISION) & MULTS_1_2(83)(PERCISION downto 1));

			MULTS_2_2(0)<=signed(MULTS_1_3(0)(PERCISION) & MULTS_1_3(0)(PERCISION downto 1))+signed(MULTS_1_4(0)(PERCISION) & MULTS_1_4(0)(PERCISION downto 1));
			MULTS_2_2(1)<=signed(MULTS_1_3(1)(PERCISION) & MULTS_1_3(1)(PERCISION downto 1))+signed(MULTS_1_4(1)(PERCISION) & MULTS_1_4(1)(PERCISION downto 1));
			MULTS_2_2(2)<=signed(MULTS_1_3(2)(PERCISION) & MULTS_1_3(2)(PERCISION downto 1))+signed(MULTS_1_4(2)(PERCISION) & MULTS_1_4(2)(PERCISION downto 1));
			MULTS_2_2(3)<=signed(MULTS_1_3(3)(PERCISION) & MULTS_1_3(3)(PERCISION downto 1))+signed(MULTS_1_4(3)(PERCISION) & MULTS_1_4(3)(PERCISION downto 1));
			MULTS_2_2(4)<=signed(MULTS_1_3(4)(PERCISION) & MULTS_1_3(4)(PERCISION downto 1))+signed(MULTS_1_4(4)(PERCISION) & MULTS_1_4(4)(PERCISION downto 1));
			MULTS_2_2(5)<=signed(MULTS_1_3(5)(PERCISION) & MULTS_1_3(5)(PERCISION downto 1))+signed(MULTS_1_4(5)(PERCISION) & MULTS_1_4(5)(PERCISION downto 1));
			MULTS_2_2(6)<=signed(MULTS_1_3(6)(PERCISION) & MULTS_1_3(6)(PERCISION downto 1))+signed(MULTS_1_4(6)(PERCISION) & MULTS_1_4(6)(PERCISION downto 1));
			MULTS_2_2(7)<=signed(MULTS_1_3(7)(PERCISION) & MULTS_1_3(7)(PERCISION downto 1))+signed(MULTS_1_4(7)(PERCISION) & MULTS_1_4(7)(PERCISION downto 1));
			MULTS_2_2(8)<=signed(MULTS_1_3(8)(PERCISION) & MULTS_1_3(8)(PERCISION downto 1))+signed(MULTS_1_4(8)(PERCISION) & MULTS_1_4(8)(PERCISION downto 1));
			MULTS_2_2(9)<=signed(MULTS_1_3(9)(PERCISION) & MULTS_1_3(9)(PERCISION downto 1))+signed(MULTS_1_4(9)(PERCISION) & MULTS_1_4(9)(PERCISION downto 1));
			MULTS_2_2(10)<=signed(MULTS_1_3(10)(PERCISION) & MULTS_1_3(10)(PERCISION downto 1))+signed(MULTS_1_4(10)(PERCISION) & MULTS_1_4(10)(PERCISION downto 1));
			MULTS_2_2(11)<=signed(MULTS_1_3(11)(PERCISION) & MULTS_1_3(11)(PERCISION downto 1))+signed(MULTS_1_4(11)(PERCISION) & MULTS_1_4(11)(PERCISION downto 1));
			MULTS_2_2(12)<=signed(MULTS_1_3(12)(PERCISION) & MULTS_1_3(12)(PERCISION downto 1))+signed(MULTS_1_4(12)(PERCISION) & MULTS_1_4(12)(PERCISION downto 1));
			MULTS_2_2(13)<=signed(MULTS_1_3(13)(PERCISION) & MULTS_1_3(13)(PERCISION downto 1))+signed(MULTS_1_4(13)(PERCISION) & MULTS_1_4(13)(PERCISION downto 1));
			MULTS_2_2(14)<=signed(MULTS_1_3(14)(PERCISION) & MULTS_1_3(14)(PERCISION downto 1))+signed(MULTS_1_4(14)(PERCISION) & MULTS_1_4(14)(PERCISION downto 1));
			MULTS_2_2(15)<=signed(MULTS_1_3(15)(PERCISION) & MULTS_1_3(15)(PERCISION downto 1))+signed(MULTS_1_4(15)(PERCISION) & MULTS_1_4(15)(PERCISION downto 1));
			MULTS_2_2(16)<=signed(MULTS_1_3(16)(PERCISION) & MULTS_1_3(16)(PERCISION downto 1))+signed(MULTS_1_4(16)(PERCISION) & MULTS_1_4(16)(PERCISION downto 1));
			MULTS_2_2(17)<=signed(MULTS_1_3(17)(PERCISION) & MULTS_1_3(17)(PERCISION downto 1))+signed(MULTS_1_4(17)(PERCISION) & MULTS_1_4(17)(PERCISION downto 1));
			MULTS_2_2(18)<=signed(MULTS_1_3(18)(PERCISION) & MULTS_1_3(18)(PERCISION downto 1))+signed(MULTS_1_4(18)(PERCISION) & MULTS_1_4(18)(PERCISION downto 1));
			MULTS_2_2(19)<=signed(MULTS_1_3(19)(PERCISION) & MULTS_1_3(19)(PERCISION downto 1))+signed(MULTS_1_4(19)(PERCISION) & MULTS_1_4(19)(PERCISION downto 1));
			MULTS_2_2(20)<=signed(MULTS_1_3(20)(PERCISION) & MULTS_1_3(20)(PERCISION downto 1))+signed(MULTS_1_4(20)(PERCISION) & MULTS_1_4(20)(PERCISION downto 1));
			MULTS_2_2(21)<=signed(MULTS_1_3(21)(PERCISION) & MULTS_1_3(21)(PERCISION downto 1))+signed(MULTS_1_4(21)(PERCISION) & MULTS_1_4(21)(PERCISION downto 1));
			MULTS_2_2(22)<=signed(MULTS_1_3(22)(PERCISION) & MULTS_1_3(22)(PERCISION downto 1))+signed(MULTS_1_4(22)(PERCISION) & MULTS_1_4(22)(PERCISION downto 1));
			MULTS_2_2(23)<=signed(MULTS_1_3(23)(PERCISION) & MULTS_1_3(23)(PERCISION downto 1))+signed(MULTS_1_4(23)(PERCISION) & MULTS_1_4(23)(PERCISION downto 1));
			MULTS_2_2(24)<=signed(MULTS_1_3(24)(PERCISION) & MULTS_1_3(24)(PERCISION downto 1))+signed(MULTS_1_4(24)(PERCISION) & MULTS_1_4(24)(PERCISION downto 1));
			MULTS_2_2(25)<=signed(MULTS_1_3(25)(PERCISION) & MULTS_1_3(25)(PERCISION downto 1))+signed(MULTS_1_4(25)(PERCISION) & MULTS_1_4(25)(PERCISION downto 1));
			MULTS_2_2(26)<=signed(MULTS_1_3(26)(PERCISION) & MULTS_1_3(26)(PERCISION downto 1))+signed(MULTS_1_4(26)(PERCISION) & MULTS_1_4(26)(PERCISION downto 1));
			MULTS_2_2(27)<=signed(MULTS_1_3(27)(PERCISION) & MULTS_1_3(27)(PERCISION downto 1))+signed(MULTS_1_4(27)(PERCISION) & MULTS_1_4(27)(PERCISION downto 1));
			MULTS_2_2(28)<=signed(MULTS_1_3(28)(PERCISION) & MULTS_1_3(28)(PERCISION downto 1))+signed(MULTS_1_4(28)(PERCISION) & MULTS_1_4(28)(PERCISION downto 1));
			MULTS_2_2(29)<=signed(MULTS_1_3(29)(PERCISION) & MULTS_1_3(29)(PERCISION downto 1))+signed(MULTS_1_4(29)(PERCISION) & MULTS_1_4(29)(PERCISION downto 1));
			MULTS_2_2(30)<=signed(MULTS_1_3(30)(PERCISION) & MULTS_1_3(30)(PERCISION downto 1))+signed(MULTS_1_4(30)(PERCISION) & MULTS_1_4(30)(PERCISION downto 1));
			MULTS_2_2(31)<=signed(MULTS_1_3(31)(PERCISION) & MULTS_1_3(31)(PERCISION downto 1))+signed(MULTS_1_4(31)(PERCISION) & MULTS_1_4(31)(PERCISION downto 1));
			MULTS_2_2(32)<=signed(MULTS_1_3(32)(PERCISION) & MULTS_1_3(32)(PERCISION downto 1))+signed(MULTS_1_4(32)(PERCISION) & MULTS_1_4(32)(PERCISION downto 1));
			MULTS_2_2(33)<=signed(MULTS_1_3(33)(PERCISION) & MULTS_1_3(33)(PERCISION downto 1))+signed(MULTS_1_4(33)(PERCISION) & MULTS_1_4(33)(PERCISION downto 1));
			MULTS_2_2(34)<=signed(MULTS_1_3(34)(PERCISION) & MULTS_1_3(34)(PERCISION downto 1))+signed(MULTS_1_4(34)(PERCISION) & MULTS_1_4(34)(PERCISION downto 1));
			MULTS_2_2(35)<=signed(MULTS_1_3(35)(PERCISION) & MULTS_1_3(35)(PERCISION downto 1))+signed(MULTS_1_4(35)(PERCISION) & MULTS_1_4(35)(PERCISION downto 1));
			MULTS_2_2(36)<=signed(MULTS_1_3(36)(PERCISION) & MULTS_1_3(36)(PERCISION downto 1))+signed(MULTS_1_4(36)(PERCISION) & MULTS_1_4(36)(PERCISION downto 1));
			MULTS_2_2(37)<=signed(MULTS_1_3(37)(PERCISION) & MULTS_1_3(37)(PERCISION downto 1))+signed(MULTS_1_4(37)(PERCISION) & MULTS_1_4(37)(PERCISION downto 1));
			MULTS_2_2(38)<=signed(MULTS_1_3(38)(PERCISION) & MULTS_1_3(38)(PERCISION downto 1))+signed(MULTS_1_4(38)(PERCISION) & MULTS_1_4(38)(PERCISION downto 1));
			MULTS_2_2(39)<=signed(MULTS_1_3(39)(PERCISION) & MULTS_1_3(39)(PERCISION downto 1))+signed(MULTS_1_4(39)(PERCISION) & MULTS_1_4(39)(PERCISION downto 1));
			MULTS_2_2(40)<=signed(MULTS_1_3(40)(PERCISION) & MULTS_1_3(40)(PERCISION downto 1))+signed(MULTS_1_4(40)(PERCISION) & MULTS_1_4(40)(PERCISION downto 1));
			MULTS_2_2(41)<=signed(MULTS_1_3(41)(PERCISION) & MULTS_1_3(41)(PERCISION downto 1))+signed(MULTS_1_4(41)(PERCISION) & MULTS_1_4(41)(PERCISION downto 1));
			MULTS_2_2(42)<=signed(MULTS_1_3(42)(PERCISION) & MULTS_1_3(42)(PERCISION downto 1))+signed(MULTS_1_4(42)(PERCISION) & MULTS_1_4(42)(PERCISION downto 1));
			MULTS_2_2(43)<=signed(MULTS_1_3(43)(PERCISION) & MULTS_1_3(43)(PERCISION downto 1))+signed(MULTS_1_4(43)(PERCISION) & MULTS_1_4(43)(PERCISION downto 1));
			MULTS_2_2(44)<=signed(MULTS_1_3(44)(PERCISION) & MULTS_1_3(44)(PERCISION downto 1))+signed(MULTS_1_4(44)(PERCISION) & MULTS_1_4(44)(PERCISION downto 1));
			MULTS_2_2(45)<=signed(MULTS_1_3(45)(PERCISION) & MULTS_1_3(45)(PERCISION downto 1))+signed(MULTS_1_4(45)(PERCISION) & MULTS_1_4(45)(PERCISION downto 1));
			MULTS_2_2(46)<=signed(MULTS_1_3(46)(PERCISION) & MULTS_1_3(46)(PERCISION downto 1))+signed(MULTS_1_4(46)(PERCISION) & MULTS_1_4(46)(PERCISION downto 1));
			MULTS_2_2(47)<=signed(MULTS_1_3(47)(PERCISION) & MULTS_1_3(47)(PERCISION downto 1))+signed(MULTS_1_4(47)(PERCISION) & MULTS_1_4(47)(PERCISION downto 1));
			MULTS_2_2(48)<=signed(MULTS_1_3(48)(PERCISION) & MULTS_1_3(48)(PERCISION downto 1))+signed(MULTS_1_4(48)(PERCISION) & MULTS_1_4(48)(PERCISION downto 1));
			MULTS_2_2(49)<=signed(MULTS_1_3(49)(PERCISION) & MULTS_1_3(49)(PERCISION downto 1))+signed(MULTS_1_4(49)(PERCISION) & MULTS_1_4(49)(PERCISION downto 1));
			MULTS_2_2(50)<=signed(MULTS_1_3(50)(PERCISION) & MULTS_1_3(50)(PERCISION downto 1))+signed(MULTS_1_4(50)(PERCISION) & MULTS_1_4(50)(PERCISION downto 1));
			MULTS_2_2(51)<=signed(MULTS_1_3(51)(PERCISION) & MULTS_1_3(51)(PERCISION downto 1))+signed(MULTS_1_4(51)(PERCISION) & MULTS_1_4(51)(PERCISION downto 1));
			MULTS_2_2(52)<=signed(MULTS_1_3(52)(PERCISION) & MULTS_1_3(52)(PERCISION downto 1))+signed(MULTS_1_4(52)(PERCISION) & MULTS_1_4(52)(PERCISION downto 1));
			MULTS_2_2(53)<=signed(MULTS_1_3(53)(PERCISION) & MULTS_1_3(53)(PERCISION downto 1))+signed(MULTS_1_4(53)(PERCISION) & MULTS_1_4(53)(PERCISION downto 1));
			MULTS_2_2(54)<=signed(MULTS_1_3(54)(PERCISION) & MULTS_1_3(54)(PERCISION downto 1))+signed(MULTS_1_4(54)(PERCISION) & MULTS_1_4(54)(PERCISION downto 1));
			MULTS_2_2(55)<=signed(MULTS_1_3(55)(PERCISION) & MULTS_1_3(55)(PERCISION downto 1))+signed(MULTS_1_4(55)(PERCISION) & MULTS_1_4(55)(PERCISION downto 1));
			MULTS_2_2(56)<=signed(MULTS_1_3(56)(PERCISION) & MULTS_1_3(56)(PERCISION downto 1))+signed(MULTS_1_4(56)(PERCISION) & MULTS_1_4(56)(PERCISION downto 1));
			MULTS_2_2(57)<=signed(MULTS_1_3(57)(PERCISION) & MULTS_1_3(57)(PERCISION downto 1))+signed(MULTS_1_4(57)(PERCISION) & MULTS_1_4(57)(PERCISION downto 1));
			MULTS_2_2(58)<=signed(MULTS_1_3(58)(PERCISION) & MULTS_1_3(58)(PERCISION downto 1))+signed(MULTS_1_4(58)(PERCISION) & MULTS_1_4(58)(PERCISION downto 1));
			MULTS_2_2(59)<=signed(MULTS_1_3(59)(PERCISION) & MULTS_1_3(59)(PERCISION downto 1))+signed(MULTS_1_4(59)(PERCISION) & MULTS_1_4(59)(PERCISION downto 1));
			MULTS_2_2(60)<=signed(MULTS_1_3(60)(PERCISION) & MULTS_1_3(60)(PERCISION downto 1))+signed(MULTS_1_4(60)(PERCISION) & MULTS_1_4(60)(PERCISION downto 1));
			MULTS_2_2(61)<=signed(MULTS_1_3(61)(PERCISION) & MULTS_1_3(61)(PERCISION downto 1))+signed(MULTS_1_4(61)(PERCISION) & MULTS_1_4(61)(PERCISION downto 1));
			MULTS_2_2(62)<=signed(MULTS_1_3(62)(PERCISION) & MULTS_1_3(62)(PERCISION downto 1))+signed(MULTS_1_4(62)(PERCISION) & MULTS_1_4(62)(PERCISION downto 1));
			MULTS_2_2(63)<=signed(MULTS_1_3(63)(PERCISION) & MULTS_1_3(63)(PERCISION downto 1))+signed(MULTS_1_4(63)(PERCISION) & MULTS_1_4(63)(PERCISION downto 1));
			MULTS_2_2(64)<=signed(MULTS_1_3(64)(PERCISION) & MULTS_1_3(64)(PERCISION downto 1))+signed(MULTS_1_4(64)(PERCISION) & MULTS_1_4(64)(PERCISION downto 1));
			MULTS_2_2(65)<=signed(MULTS_1_3(65)(PERCISION) & MULTS_1_3(65)(PERCISION downto 1))+signed(MULTS_1_4(65)(PERCISION) & MULTS_1_4(65)(PERCISION downto 1));
			MULTS_2_2(66)<=signed(MULTS_1_3(66)(PERCISION) & MULTS_1_3(66)(PERCISION downto 1))+signed(MULTS_1_4(66)(PERCISION) & MULTS_1_4(66)(PERCISION downto 1));
			MULTS_2_2(67)<=signed(MULTS_1_3(67)(PERCISION) & MULTS_1_3(67)(PERCISION downto 1))+signed(MULTS_1_4(67)(PERCISION) & MULTS_1_4(67)(PERCISION downto 1));
			MULTS_2_2(68)<=signed(MULTS_1_3(68)(PERCISION) & MULTS_1_3(68)(PERCISION downto 1))+signed(MULTS_1_4(68)(PERCISION) & MULTS_1_4(68)(PERCISION downto 1));
			MULTS_2_2(69)<=signed(MULTS_1_3(69)(PERCISION) & MULTS_1_3(69)(PERCISION downto 1))+signed(MULTS_1_4(69)(PERCISION) & MULTS_1_4(69)(PERCISION downto 1));
			MULTS_2_2(70)<=signed(MULTS_1_3(70)(PERCISION) & MULTS_1_3(70)(PERCISION downto 1))+signed(MULTS_1_4(70)(PERCISION) & MULTS_1_4(70)(PERCISION downto 1));
			MULTS_2_2(71)<=signed(MULTS_1_3(71)(PERCISION) & MULTS_1_3(71)(PERCISION downto 1))+signed(MULTS_1_4(71)(PERCISION) & MULTS_1_4(71)(PERCISION downto 1));
			MULTS_2_2(72)<=signed(MULTS_1_3(72)(PERCISION) & MULTS_1_3(72)(PERCISION downto 1))+signed(MULTS_1_4(72)(PERCISION) & MULTS_1_4(72)(PERCISION downto 1));
			MULTS_2_2(73)<=signed(MULTS_1_3(73)(PERCISION) & MULTS_1_3(73)(PERCISION downto 1))+signed(MULTS_1_4(73)(PERCISION) & MULTS_1_4(73)(PERCISION downto 1));
			MULTS_2_2(74)<=signed(MULTS_1_3(74)(PERCISION) & MULTS_1_3(74)(PERCISION downto 1))+signed(MULTS_1_4(74)(PERCISION) & MULTS_1_4(74)(PERCISION downto 1));
			MULTS_2_2(75)<=signed(MULTS_1_3(75)(PERCISION) & MULTS_1_3(75)(PERCISION downto 1))+signed(MULTS_1_4(75)(PERCISION) & MULTS_1_4(75)(PERCISION downto 1));
			MULTS_2_2(76)<=signed(MULTS_1_3(76)(PERCISION) & MULTS_1_3(76)(PERCISION downto 1))+signed(MULTS_1_4(76)(PERCISION) & MULTS_1_4(76)(PERCISION downto 1));
			MULTS_2_2(77)<=signed(MULTS_1_3(77)(PERCISION) & MULTS_1_3(77)(PERCISION downto 1))+signed(MULTS_1_4(77)(PERCISION) & MULTS_1_4(77)(PERCISION downto 1));
			MULTS_2_2(78)<=signed(MULTS_1_3(78)(PERCISION) & MULTS_1_3(78)(PERCISION downto 1))+signed(MULTS_1_4(78)(PERCISION) & MULTS_1_4(78)(PERCISION downto 1));
			MULTS_2_2(79)<=signed(MULTS_1_3(79)(PERCISION) & MULTS_1_3(79)(PERCISION downto 1))+signed(MULTS_1_4(79)(PERCISION) & MULTS_1_4(79)(PERCISION downto 1));
			MULTS_2_2(80)<=signed(MULTS_1_3(80)(PERCISION) & MULTS_1_3(80)(PERCISION downto 1))+signed(MULTS_1_4(80)(PERCISION) & MULTS_1_4(80)(PERCISION downto 1));
			MULTS_2_2(81)<=signed(MULTS_1_3(81)(PERCISION) & MULTS_1_3(81)(PERCISION downto 1))+signed(MULTS_1_4(81)(PERCISION) & MULTS_1_4(81)(PERCISION downto 1));
			MULTS_2_2(82)<=signed(MULTS_1_3(82)(PERCISION) & MULTS_1_3(82)(PERCISION downto 1))+signed(MULTS_1_4(82)(PERCISION) & MULTS_1_4(82)(PERCISION downto 1));
			MULTS_2_2(83)<=signed(MULTS_1_3(83)(PERCISION) & MULTS_1_3(83)(PERCISION downto 1))+signed(MULTS_1_4(83)(PERCISION) & MULTS_1_4(83)(PERCISION downto 1));

			MULTS_2_3(0)<=signed(MULTS_1_5(0)(PERCISION) & MULTS_1_5(0)(PERCISION downto 1))+signed(MULTS_1_6(0)(PERCISION) & MULTS_1_6(0)(PERCISION downto 1));
			MULTS_2_3(1)<=signed(MULTS_1_5(1)(PERCISION) & MULTS_1_5(1)(PERCISION downto 1))+signed(MULTS_1_6(1)(PERCISION) & MULTS_1_6(1)(PERCISION downto 1));
			MULTS_2_3(2)<=signed(MULTS_1_5(2)(PERCISION) & MULTS_1_5(2)(PERCISION downto 1))+signed(MULTS_1_6(2)(PERCISION) & MULTS_1_6(2)(PERCISION downto 1));
			MULTS_2_3(3)<=signed(MULTS_1_5(3)(PERCISION) & MULTS_1_5(3)(PERCISION downto 1))+signed(MULTS_1_6(3)(PERCISION) & MULTS_1_6(3)(PERCISION downto 1));
			MULTS_2_3(4)<=signed(MULTS_1_5(4)(PERCISION) & MULTS_1_5(4)(PERCISION downto 1))+signed(MULTS_1_6(4)(PERCISION) & MULTS_1_6(4)(PERCISION downto 1));
			MULTS_2_3(5)<=signed(MULTS_1_5(5)(PERCISION) & MULTS_1_5(5)(PERCISION downto 1))+signed(MULTS_1_6(5)(PERCISION) & MULTS_1_6(5)(PERCISION downto 1));
			MULTS_2_3(6)<=signed(MULTS_1_5(6)(PERCISION) & MULTS_1_5(6)(PERCISION downto 1))+signed(MULTS_1_6(6)(PERCISION) & MULTS_1_6(6)(PERCISION downto 1));
			MULTS_2_3(7)<=signed(MULTS_1_5(7)(PERCISION) & MULTS_1_5(7)(PERCISION downto 1))+signed(MULTS_1_6(7)(PERCISION) & MULTS_1_6(7)(PERCISION downto 1));
			MULTS_2_3(8)<=signed(MULTS_1_5(8)(PERCISION) & MULTS_1_5(8)(PERCISION downto 1))+signed(MULTS_1_6(8)(PERCISION) & MULTS_1_6(8)(PERCISION downto 1));
			MULTS_2_3(9)<=signed(MULTS_1_5(9)(PERCISION) & MULTS_1_5(9)(PERCISION downto 1))+signed(MULTS_1_6(9)(PERCISION) & MULTS_1_6(9)(PERCISION downto 1));
			MULTS_2_3(10)<=signed(MULTS_1_5(10)(PERCISION) & MULTS_1_5(10)(PERCISION downto 1))+signed(MULTS_1_6(10)(PERCISION) & MULTS_1_6(10)(PERCISION downto 1));
			MULTS_2_3(11)<=signed(MULTS_1_5(11)(PERCISION) & MULTS_1_5(11)(PERCISION downto 1))+signed(MULTS_1_6(11)(PERCISION) & MULTS_1_6(11)(PERCISION downto 1));
			MULTS_2_3(12)<=signed(MULTS_1_5(12)(PERCISION) & MULTS_1_5(12)(PERCISION downto 1))+signed(MULTS_1_6(12)(PERCISION) & MULTS_1_6(12)(PERCISION downto 1));
			MULTS_2_3(13)<=signed(MULTS_1_5(13)(PERCISION) & MULTS_1_5(13)(PERCISION downto 1))+signed(MULTS_1_6(13)(PERCISION) & MULTS_1_6(13)(PERCISION downto 1));
			MULTS_2_3(14)<=signed(MULTS_1_5(14)(PERCISION) & MULTS_1_5(14)(PERCISION downto 1))+signed(MULTS_1_6(14)(PERCISION) & MULTS_1_6(14)(PERCISION downto 1));
			MULTS_2_3(15)<=signed(MULTS_1_5(15)(PERCISION) & MULTS_1_5(15)(PERCISION downto 1))+signed(MULTS_1_6(15)(PERCISION) & MULTS_1_6(15)(PERCISION downto 1));
			MULTS_2_3(16)<=signed(MULTS_1_5(16)(PERCISION) & MULTS_1_5(16)(PERCISION downto 1))+signed(MULTS_1_6(16)(PERCISION) & MULTS_1_6(16)(PERCISION downto 1));
			MULTS_2_3(17)<=signed(MULTS_1_5(17)(PERCISION) & MULTS_1_5(17)(PERCISION downto 1))+signed(MULTS_1_6(17)(PERCISION) & MULTS_1_6(17)(PERCISION downto 1));
			MULTS_2_3(18)<=signed(MULTS_1_5(18)(PERCISION) & MULTS_1_5(18)(PERCISION downto 1))+signed(MULTS_1_6(18)(PERCISION) & MULTS_1_6(18)(PERCISION downto 1));
			MULTS_2_3(19)<=signed(MULTS_1_5(19)(PERCISION) & MULTS_1_5(19)(PERCISION downto 1))+signed(MULTS_1_6(19)(PERCISION) & MULTS_1_6(19)(PERCISION downto 1));
			MULTS_2_3(20)<=signed(MULTS_1_5(20)(PERCISION) & MULTS_1_5(20)(PERCISION downto 1))+signed(MULTS_1_6(20)(PERCISION) & MULTS_1_6(20)(PERCISION downto 1));
			MULTS_2_3(21)<=signed(MULTS_1_5(21)(PERCISION) & MULTS_1_5(21)(PERCISION downto 1))+signed(MULTS_1_6(21)(PERCISION) & MULTS_1_6(21)(PERCISION downto 1));
			MULTS_2_3(22)<=signed(MULTS_1_5(22)(PERCISION) & MULTS_1_5(22)(PERCISION downto 1))+signed(MULTS_1_6(22)(PERCISION) & MULTS_1_6(22)(PERCISION downto 1));
			MULTS_2_3(23)<=signed(MULTS_1_5(23)(PERCISION) & MULTS_1_5(23)(PERCISION downto 1))+signed(MULTS_1_6(23)(PERCISION) & MULTS_1_6(23)(PERCISION downto 1));
			MULTS_2_3(24)<=signed(MULTS_1_5(24)(PERCISION) & MULTS_1_5(24)(PERCISION downto 1))+signed(MULTS_1_6(24)(PERCISION) & MULTS_1_6(24)(PERCISION downto 1));
			MULTS_2_3(25)<=signed(MULTS_1_5(25)(PERCISION) & MULTS_1_5(25)(PERCISION downto 1))+signed(MULTS_1_6(25)(PERCISION) & MULTS_1_6(25)(PERCISION downto 1));
			MULTS_2_3(26)<=signed(MULTS_1_5(26)(PERCISION) & MULTS_1_5(26)(PERCISION downto 1))+signed(MULTS_1_6(26)(PERCISION) & MULTS_1_6(26)(PERCISION downto 1));
			MULTS_2_3(27)<=signed(MULTS_1_5(27)(PERCISION) & MULTS_1_5(27)(PERCISION downto 1))+signed(MULTS_1_6(27)(PERCISION) & MULTS_1_6(27)(PERCISION downto 1));
			MULTS_2_3(28)<=signed(MULTS_1_5(28)(PERCISION) & MULTS_1_5(28)(PERCISION downto 1))+signed(MULTS_1_6(28)(PERCISION) & MULTS_1_6(28)(PERCISION downto 1));
			MULTS_2_3(29)<=signed(MULTS_1_5(29)(PERCISION) & MULTS_1_5(29)(PERCISION downto 1))+signed(MULTS_1_6(29)(PERCISION) & MULTS_1_6(29)(PERCISION downto 1));
			MULTS_2_3(30)<=signed(MULTS_1_5(30)(PERCISION) & MULTS_1_5(30)(PERCISION downto 1))+signed(MULTS_1_6(30)(PERCISION) & MULTS_1_6(30)(PERCISION downto 1));
			MULTS_2_3(31)<=signed(MULTS_1_5(31)(PERCISION) & MULTS_1_5(31)(PERCISION downto 1))+signed(MULTS_1_6(31)(PERCISION) & MULTS_1_6(31)(PERCISION downto 1));
			MULTS_2_3(32)<=signed(MULTS_1_5(32)(PERCISION) & MULTS_1_5(32)(PERCISION downto 1))+signed(MULTS_1_6(32)(PERCISION) & MULTS_1_6(32)(PERCISION downto 1));
			MULTS_2_3(33)<=signed(MULTS_1_5(33)(PERCISION) & MULTS_1_5(33)(PERCISION downto 1))+signed(MULTS_1_6(33)(PERCISION) & MULTS_1_6(33)(PERCISION downto 1));
			MULTS_2_3(34)<=signed(MULTS_1_5(34)(PERCISION) & MULTS_1_5(34)(PERCISION downto 1))+signed(MULTS_1_6(34)(PERCISION) & MULTS_1_6(34)(PERCISION downto 1));
			MULTS_2_3(35)<=signed(MULTS_1_5(35)(PERCISION) & MULTS_1_5(35)(PERCISION downto 1))+signed(MULTS_1_6(35)(PERCISION) & MULTS_1_6(35)(PERCISION downto 1));
			MULTS_2_3(36)<=signed(MULTS_1_5(36)(PERCISION) & MULTS_1_5(36)(PERCISION downto 1))+signed(MULTS_1_6(36)(PERCISION) & MULTS_1_6(36)(PERCISION downto 1));
			MULTS_2_3(37)<=signed(MULTS_1_5(37)(PERCISION) & MULTS_1_5(37)(PERCISION downto 1))+signed(MULTS_1_6(37)(PERCISION) & MULTS_1_6(37)(PERCISION downto 1));
			MULTS_2_3(38)<=signed(MULTS_1_5(38)(PERCISION) & MULTS_1_5(38)(PERCISION downto 1))+signed(MULTS_1_6(38)(PERCISION) & MULTS_1_6(38)(PERCISION downto 1));
			MULTS_2_3(39)<=signed(MULTS_1_5(39)(PERCISION) & MULTS_1_5(39)(PERCISION downto 1))+signed(MULTS_1_6(39)(PERCISION) & MULTS_1_6(39)(PERCISION downto 1));
			MULTS_2_3(40)<=signed(MULTS_1_5(40)(PERCISION) & MULTS_1_5(40)(PERCISION downto 1))+signed(MULTS_1_6(40)(PERCISION) & MULTS_1_6(40)(PERCISION downto 1));
			MULTS_2_3(41)<=signed(MULTS_1_5(41)(PERCISION) & MULTS_1_5(41)(PERCISION downto 1))+signed(MULTS_1_6(41)(PERCISION) & MULTS_1_6(41)(PERCISION downto 1));
			MULTS_2_3(42)<=signed(MULTS_1_5(42)(PERCISION) & MULTS_1_5(42)(PERCISION downto 1))+signed(MULTS_1_6(42)(PERCISION) & MULTS_1_6(42)(PERCISION downto 1));
			MULTS_2_3(43)<=signed(MULTS_1_5(43)(PERCISION) & MULTS_1_5(43)(PERCISION downto 1))+signed(MULTS_1_6(43)(PERCISION) & MULTS_1_6(43)(PERCISION downto 1));
			MULTS_2_3(44)<=signed(MULTS_1_5(44)(PERCISION) & MULTS_1_5(44)(PERCISION downto 1))+signed(MULTS_1_6(44)(PERCISION) & MULTS_1_6(44)(PERCISION downto 1));
			MULTS_2_3(45)<=signed(MULTS_1_5(45)(PERCISION) & MULTS_1_5(45)(PERCISION downto 1))+signed(MULTS_1_6(45)(PERCISION) & MULTS_1_6(45)(PERCISION downto 1));
			MULTS_2_3(46)<=signed(MULTS_1_5(46)(PERCISION) & MULTS_1_5(46)(PERCISION downto 1))+signed(MULTS_1_6(46)(PERCISION) & MULTS_1_6(46)(PERCISION downto 1));
			MULTS_2_3(47)<=signed(MULTS_1_5(47)(PERCISION) & MULTS_1_5(47)(PERCISION downto 1))+signed(MULTS_1_6(47)(PERCISION) & MULTS_1_6(47)(PERCISION downto 1));
			MULTS_2_3(48)<=signed(MULTS_1_5(48)(PERCISION) & MULTS_1_5(48)(PERCISION downto 1))+signed(MULTS_1_6(48)(PERCISION) & MULTS_1_6(48)(PERCISION downto 1));
			MULTS_2_3(49)<=signed(MULTS_1_5(49)(PERCISION) & MULTS_1_5(49)(PERCISION downto 1))+signed(MULTS_1_6(49)(PERCISION) & MULTS_1_6(49)(PERCISION downto 1));
			MULTS_2_3(50)<=signed(MULTS_1_5(50)(PERCISION) & MULTS_1_5(50)(PERCISION downto 1))+signed(MULTS_1_6(50)(PERCISION) & MULTS_1_6(50)(PERCISION downto 1));
			MULTS_2_3(51)<=signed(MULTS_1_5(51)(PERCISION) & MULTS_1_5(51)(PERCISION downto 1))+signed(MULTS_1_6(51)(PERCISION) & MULTS_1_6(51)(PERCISION downto 1));
			MULTS_2_3(52)<=signed(MULTS_1_5(52)(PERCISION) & MULTS_1_5(52)(PERCISION downto 1))+signed(MULTS_1_6(52)(PERCISION) & MULTS_1_6(52)(PERCISION downto 1));
			MULTS_2_3(53)<=signed(MULTS_1_5(53)(PERCISION) & MULTS_1_5(53)(PERCISION downto 1))+signed(MULTS_1_6(53)(PERCISION) & MULTS_1_6(53)(PERCISION downto 1));
			MULTS_2_3(54)<=signed(MULTS_1_5(54)(PERCISION) & MULTS_1_5(54)(PERCISION downto 1))+signed(MULTS_1_6(54)(PERCISION) & MULTS_1_6(54)(PERCISION downto 1));
			MULTS_2_3(55)<=signed(MULTS_1_5(55)(PERCISION) & MULTS_1_5(55)(PERCISION downto 1))+signed(MULTS_1_6(55)(PERCISION) & MULTS_1_6(55)(PERCISION downto 1));
			MULTS_2_3(56)<=signed(MULTS_1_5(56)(PERCISION) & MULTS_1_5(56)(PERCISION downto 1))+signed(MULTS_1_6(56)(PERCISION) & MULTS_1_6(56)(PERCISION downto 1));
			MULTS_2_3(57)<=signed(MULTS_1_5(57)(PERCISION) & MULTS_1_5(57)(PERCISION downto 1))+signed(MULTS_1_6(57)(PERCISION) & MULTS_1_6(57)(PERCISION downto 1));
			MULTS_2_3(58)<=signed(MULTS_1_5(58)(PERCISION) & MULTS_1_5(58)(PERCISION downto 1))+signed(MULTS_1_6(58)(PERCISION) & MULTS_1_6(58)(PERCISION downto 1));
			MULTS_2_3(59)<=signed(MULTS_1_5(59)(PERCISION) & MULTS_1_5(59)(PERCISION downto 1))+signed(MULTS_1_6(59)(PERCISION) & MULTS_1_6(59)(PERCISION downto 1));
			MULTS_2_3(60)<=signed(MULTS_1_5(60)(PERCISION) & MULTS_1_5(60)(PERCISION downto 1))+signed(MULTS_1_6(60)(PERCISION) & MULTS_1_6(60)(PERCISION downto 1));
			MULTS_2_3(61)<=signed(MULTS_1_5(61)(PERCISION) & MULTS_1_5(61)(PERCISION downto 1))+signed(MULTS_1_6(61)(PERCISION) & MULTS_1_6(61)(PERCISION downto 1));
			MULTS_2_3(62)<=signed(MULTS_1_5(62)(PERCISION) & MULTS_1_5(62)(PERCISION downto 1))+signed(MULTS_1_6(62)(PERCISION) & MULTS_1_6(62)(PERCISION downto 1));
			MULTS_2_3(63)<=signed(MULTS_1_5(63)(PERCISION) & MULTS_1_5(63)(PERCISION downto 1))+signed(MULTS_1_6(63)(PERCISION) & MULTS_1_6(63)(PERCISION downto 1));
			MULTS_2_3(64)<=signed(MULTS_1_5(64)(PERCISION) & MULTS_1_5(64)(PERCISION downto 1))+signed(MULTS_1_6(64)(PERCISION) & MULTS_1_6(64)(PERCISION downto 1));
			MULTS_2_3(65)<=signed(MULTS_1_5(65)(PERCISION) & MULTS_1_5(65)(PERCISION downto 1))+signed(MULTS_1_6(65)(PERCISION) & MULTS_1_6(65)(PERCISION downto 1));
			MULTS_2_3(66)<=signed(MULTS_1_5(66)(PERCISION) & MULTS_1_5(66)(PERCISION downto 1))+signed(MULTS_1_6(66)(PERCISION) & MULTS_1_6(66)(PERCISION downto 1));
			MULTS_2_3(67)<=signed(MULTS_1_5(67)(PERCISION) & MULTS_1_5(67)(PERCISION downto 1))+signed(MULTS_1_6(67)(PERCISION) & MULTS_1_6(67)(PERCISION downto 1));
			MULTS_2_3(68)<=signed(MULTS_1_5(68)(PERCISION) & MULTS_1_5(68)(PERCISION downto 1))+signed(MULTS_1_6(68)(PERCISION) & MULTS_1_6(68)(PERCISION downto 1));
			MULTS_2_3(69)<=signed(MULTS_1_5(69)(PERCISION) & MULTS_1_5(69)(PERCISION downto 1))+signed(MULTS_1_6(69)(PERCISION) & MULTS_1_6(69)(PERCISION downto 1));
			MULTS_2_3(70)<=signed(MULTS_1_5(70)(PERCISION) & MULTS_1_5(70)(PERCISION downto 1))+signed(MULTS_1_6(70)(PERCISION) & MULTS_1_6(70)(PERCISION downto 1));
			MULTS_2_3(71)<=signed(MULTS_1_5(71)(PERCISION) & MULTS_1_5(71)(PERCISION downto 1))+signed(MULTS_1_6(71)(PERCISION) & MULTS_1_6(71)(PERCISION downto 1));
			MULTS_2_3(72)<=signed(MULTS_1_5(72)(PERCISION) & MULTS_1_5(72)(PERCISION downto 1))+signed(MULTS_1_6(72)(PERCISION) & MULTS_1_6(72)(PERCISION downto 1));
			MULTS_2_3(73)<=signed(MULTS_1_5(73)(PERCISION) & MULTS_1_5(73)(PERCISION downto 1))+signed(MULTS_1_6(73)(PERCISION) & MULTS_1_6(73)(PERCISION downto 1));
			MULTS_2_3(74)<=signed(MULTS_1_5(74)(PERCISION) & MULTS_1_5(74)(PERCISION downto 1))+signed(MULTS_1_6(74)(PERCISION) & MULTS_1_6(74)(PERCISION downto 1));
			MULTS_2_3(75)<=signed(MULTS_1_5(75)(PERCISION) & MULTS_1_5(75)(PERCISION downto 1))+signed(MULTS_1_6(75)(PERCISION) & MULTS_1_6(75)(PERCISION downto 1));
			MULTS_2_3(76)<=signed(MULTS_1_5(76)(PERCISION) & MULTS_1_5(76)(PERCISION downto 1))+signed(MULTS_1_6(76)(PERCISION) & MULTS_1_6(76)(PERCISION downto 1));
			MULTS_2_3(77)<=signed(MULTS_1_5(77)(PERCISION) & MULTS_1_5(77)(PERCISION downto 1))+signed(MULTS_1_6(77)(PERCISION) & MULTS_1_6(77)(PERCISION downto 1));
			MULTS_2_3(78)<=signed(MULTS_1_5(78)(PERCISION) & MULTS_1_5(78)(PERCISION downto 1))+signed(MULTS_1_6(78)(PERCISION) & MULTS_1_6(78)(PERCISION downto 1));
			MULTS_2_3(79)<=signed(MULTS_1_5(79)(PERCISION) & MULTS_1_5(79)(PERCISION downto 1))+signed(MULTS_1_6(79)(PERCISION) & MULTS_1_6(79)(PERCISION downto 1));
			MULTS_2_3(80)<=signed(MULTS_1_5(80)(PERCISION) & MULTS_1_5(80)(PERCISION downto 1))+signed(MULTS_1_6(80)(PERCISION) & MULTS_1_6(80)(PERCISION downto 1));
			MULTS_2_3(81)<=signed(MULTS_1_5(81)(PERCISION) & MULTS_1_5(81)(PERCISION downto 1))+signed(MULTS_1_6(81)(PERCISION) & MULTS_1_6(81)(PERCISION downto 1));
			MULTS_2_3(82)<=signed(MULTS_1_5(82)(PERCISION) & MULTS_1_5(82)(PERCISION downto 1))+signed(MULTS_1_6(82)(PERCISION) & MULTS_1_6(82)(PERCISION downto 1));
			MULTS_2_3(83)<=signed(MULTS_1_5(83)(PERCISION) & MULTS_1_5(83)(PERCISION downto 1))+signed(MULTS_1_6(83)(PERCISION) & MULTS_1_6(83)(PERCISION downto 1));

			MULTS_2_4(0)<=signed(MULTS_1_7(0)(PERCISION) & MULTS_1_7(0)(PERCISION downto 1))+signed(MULTS_1_8(0)(PERCISION) & MULTS_1_8(0)(PERCISION downto 1));
			MULTS_2_4(1)<=signed(MULTS_1_7(1)(PERCISION) & MULTS_1_7(1)(PERCISION downto 1))+signed(MULTS_1_8(1)(PERCISION) & MULTS_1_8(1)(PERCISION downto 1));
			MULTS_2_4(2)<=signed(MULTS_1_7(2)(PERCISION) & MULTS_1_7(2)(PERCISION downto 1))+signed(MULTS_1_8(2)(PERCISION) & MULTS_1_8(2)(PERCISION downto 1));
			MULTS_2_4(3)<=signed(MULTS_1_7(3)(PERCISION) & MULTS_1_7(3)(PERCISION downto 1))+signed(MULTS_1_8(3)(PERCISION) & MULTS_1_8(3)(PERCISION downto 1));
			MULTS_2_4(4)<=signed(MULTS_1_7(4)(PERCISION) & MULTS_1_7(4)(PERCISION downto 1))+signed(MULTS_1_8(4)(PERCISION) & MULTS_1_8(4)(PERCISION downto 1));
			MULTS_2_4(5)<=signed(MULTS_1_7(5)(PERCISION) & MULTS_1_7(5)(PERCISION downto 1))+signed(MULTS_1_8(5)(PERCISION) & MULTS_1_8(5)(PERCISION downto 1));
			MULTS_2_4(6)<=signed(MULTS_1_7(6)(PERCISION) & MULTS_1_7(6)(PERCISION downto 1))+signed(MULTS_1_8(6)(PERCISION) & MULTS_1_8(6)(PERCISION downto 1));
			MULTS_2_4(7)<=signed(MULTS_1_7(7)(PERCISION) & MULTS_1_7(7)(PERCISION downto 1))+signed(MULTS_1_8(7)(PERCISION) & MULTS_1_8(7)(PERCISION downto 1));
			MULTS_2_4(8)<=signed(MULTS_1_7(8)(PERCISION) & MULTS_1_7(8)(PERCISION downto 1))+signed(MULTS_1_8(8)(PERCISION) & MULTS_1_8(8)(PERCISION downto 1));
			MULTS_2_4(9)<=signed(MULTS_1_7(9)(PERCISION) & MULTS_1_7(9)(PERCISION downto 1))+signed(MULTS_1_8(9)(PERCISION) & MULTS_1_8(9)(PERCISION downto 1));
			MULTS_2_4(10)<=signed(MULTS_1_7(10)(PERCISION) & MULTS_1_7(10)(PERCISION downto 1))+signed(MULTS_1_8(10)(PERCISION) & MULTS_1_8(10)(PERCISION downto 1));
			MULTS_2_4(11)<=signed(MULTS_1_7(11)(PERCISION) & MULTS_1_7(11)(PERCISION downto 1))+signed(MULTS_1_8(11)(PERCISION) & MULTS_1_8(11)(PERCISION downto 1));
			MULTS_2_4(12)<=signed(MULTS_1_7(12)(PERCISION) & MULTS_1_7(12)(PERCISION downto 1))+signed(MULTS_1_8(12)(PERCISION) & MULTS_1_8(12)(PERCISION downto 1));
			MULTS_2_4(13)<=signed(MULTS_1_7(13)(PERCISION) & MULTS_1_7(13)(PERCISION downto 1))+signed(MULTS_1_8(13)(PERCISION) & MULTS_1_8(13)(PERCISION downto 1));
			MULTS_2_4(14)<=signed(MULTS_1_7(14)(PERCISION) & MULTS_1_7(14)(PERCISION downto 1))+signed(MULTS_1_8(14)(PERCISION) & MULTS_1_8(14)(PERCISION downto 1));
			MULTS_2_4(15)<=signed(MULTS_1_7(15)(PERCISION) & MULTS_1_7(15)(PERCISION downto 1))+signed(MULTS_1_8(15)(PERCISION) & MULTS_1_8(15)(PERCISION downto 1));
			MULTS_2_4(16)<=signed(MULTS_1_7(16)(PERCISION) & MULTS_1_7(16)(PERCISION downto 1))+signed(MULTS_1_8(16)(PERCISION) & MULTS_1_8(16)(PERCISION downto 1));
			MULTS_2_4(17)<=signed(MULTS_1_7(17)(PERCISION) & MULTS_1_7(17)(PERCISION downto 1))+signed(MULTS_1_8(17)(PERCISION) & MULTS_1_8(17)(PERCISION downto 1));
			MULTS_2_4(18)<=signed(MULTS_1_7(18)(PERCISION) & MULTS_1_7(18)(PERCISION downto 1))+signed(MULTS_1_8(18)(PERCISION) & MULTS_1_8(18)(PERCISION downto 1));
			MULTS_2_4(19)<=signed(MULTS_1_7(19)(PERCISION) & MULTS_1_7(19)(PERCISION downto 1))+signed(MULTS_1_8(19)(PERCISION) & MULTS_1_8(19)(PERCISION downto 1));
			MULTS_2_4(20)<=signed(MULTS_1_7(20)(PERCISION) & MULTS_1_7(20)(PERCISION downto 1))+signed(MULTS_1_8(20)(PERCISION) & MULTS_1_8(20)(PERCISION downto 1));
			MULTS_2_4(21)<=signed(MULTS_1_7(21)(PERCISION) & MULTS_1_7(21)(PERCISION downto 1))+signed(MULTS_1_8(21)(PERCISION) & MULTS_1_8(21)(PERCISION downto 1));
			MULTS_2_4(22)<=signed(MULTS_1_7(22)(PERCISION) & MULTS_1_7(22)(PERCISION downto 1))+signed(MULTS_1_8(22)(PERCISION) & MULTS_1_8(22)(PERCISION downto 1));
			MULTS_2_4(23)<=signed(MULTS_1_7(23)(PERCISION) & MULTS_1_7(23)(PERCISION downto 1))+signed(MULTS_1_8(23)(PERCISION) & MULTS_1_8(23)(PERCISION downto 1));
			MULTS_2_4(24)<=signed(MULTS_1_7(24)(PERCISION) & MULTS_1_7(24)(PERCISION downto 1))+signed(MULTS_1_8(24)(PERCISION) & MULTS_1_8(24)(PERCISION downto 1));
			MULTS_2_4(25)<=signed(MULTS_1_7(25)(PERCISION) & MULTS_1_7(25)(PERCISION downto 1))+signed(MULTS_1_8(25)(PERCISION) & MULTS_1_8(25)(PERCISION downto 1));
			MULTS_2_4(26)<=signed(MULTS_1_7(26)(PERCISION) & MULTS_1_7(26)(PERCISION downto 1))+signed(MULTS_1_8(26)(PERCISION) & MULTS_1_8(26)(PERCISION downto 1));
			MULTS_2_4(27)<=signed(MULTS_1_7(27)(PERCISION) & MULTS_1_7(27)(PERCISION downto 1))+signed(MULTS_1_8(27)(PERCISION) & MULTS_1_8(27)(PERCISION downto 1));
			MULTS_2_4(28)<=signed(MULTS_1_7(28)(PERCISION) & MULTS_1_7(28)(PERCISION downto 1))+signed(MULTS_1_8(28)(PERCISION) & MULTS_1_8(28)(PERCISION downto 1));
			MULTS_2_4(29)<=signed(MULTS_1_7(29)(PERCISION) & MULTS_1_7(29)(PERCISION downto 1))+signed(MULTS_1_8(29)(PERCISION) & MULTS_1_8(29)(PERCISION downto 1));
			MULTS_2_4(30)<=signed(MULTS_1_7(30)(PERCISION) & MULTS_1_7(30)(PERCISION downto 1))+signed(MULTS_1_8(30)(PERCISION) & MULTS_1_8(30)(PERCISION downto 1));
			MULTS_2_4(31)<=signed(MULTS_1_7(31)(PERCISION) & MULTS_1_7(31)(PERCISION downto 1))+signed(MULTS_1_8(31)(PERCISION) & MULTS_1_8(31)(PERCISION downto 1));
			MULTS_2_4(32)<=signed(MULTS_1_7(32)(PERCISION) & MULTS_1_7(32)(PERCISION downto 1))+signed(MULTS_1_8(32)(PERCISION) & MULTS_1_8(32)(PERCISION downto 1));
			MULTS_2_4(33)<=signed(MULTS_1_7(33)(PERCISION) & MULTS_1_7(33)(PERCISION downto 1))+signed(MULTS_1_8(33)(PERCISION) & MULTS_1_8(33)(PERCISION downto 1));
			MULTS_2_4(34)<=signed(MULTS_1_7(34)(PERCISION) & MULTS_1_7(34)(PERCISION downto 1))+signed(MULTS_1_8(34)(PERCISION) & MULTS_1_8(34)(PERCISION downto 1));
			MULTS_2_4(35)<=signed(MULTS_1_7(35)(PERCISION) & MULTS_1_7(35)(PERCISION downto 1))+signed(MULTS_1_8(35)(PERCISION) & MULTS_1_8(35)(PERCISION downto 1));
			MULTS_2_4(36)<=signed(MULTS_1_7(36)(PERCISION) & MULTS_1_7(36)(PERCISION downto 1))+signed(MULTS_1_8(36)(PERCISION) & MULTS_1_8(36)(PERCISION downto 1));
			MULTS_2_4(37)<=signed(MULTS_1_7(37)(PERCISION) & MULTS_1_7(37)(PERCISION downto 1))+signed(MULTS_1_8(37)(PERCISION) & MULTS_1_8(37)(PERCISION downto 1));
			MULTS_2_4(38)<=signed(MULTS_1_7(38)(PERCISION) & MULTS_1_7(38)(PERCISION downto 1))+signed(MULTS_1_8(38)(PERCISION) & MULTS_1_8(38)(PERCISION downto 1));
			MULTS_2_4(39)<=signed(MULTS_1_7(39)(PERCISION) & MULTS_1_7(39)(PERCISION downto 1))+signed(MULTS_1_8(39)(PERCISION) & MULTS_1_8(39)(PERCISION downto 1));
			MULTS_2_4(40)<=signed(MULTS_1_7(40)(PERCISION) & MULTS_1_7(40)(PERCISION downto 1))+signed(MULTS_1_8(40)(PERCISION) & MULTS_1_8(40)(PERCISION downto 1));
			MULTS_2_4(41)<=signed(MULTS_1_7(41)(PERCISION) & MULTS_1_7(41)(PERCISION downto 1))+signed(MULTS_1_8(41)(PERCISION) & MULTS_1_8(41)(PERCISION downto 1));
			MULTS_2_4(42)<=signed(MULTS_1_7(42)(PERCISION) & MULTS_1_7(42)(PERCISION downto 1))+signed(MULTS_1_8(42)(PERCISION) & MULTS_1_8(42)(PERCISION downto 1));
			MULTS_2_4(43)<=signed(MULTS_1_7(43)(PERCISION) & MULTS_1_7(43)(PERCISION downto 1))+signed(MULTS_1_8(43)(PERCISION) & MULTS_1_8(43)(PERCISION downto 1));
			MULTS_2_4(44)<=signed(MULTS_1_7(44)(PERCISION) & MULTS_1_7(44)(PERCISION downto 1))+signed(MULTS_1_8(44)(PERCISION) & MULTS_1_8(44)(PERCISION downto 1));
			MULTS_2_4(45)<=signed(MULTS_1_7(45)(PERCISION) & MULTS_1_7(45)(PERCISION downto 1))+signed(MULTS_1_8(45)(PERCISION) & MULTS_1_8(45)(PERCISION downto 1));
			MULTS_2_4(46)<=signed(MULTS_1_7(46)(PERCISION) & MULTS_1_7(46)(PERCISION downto 1))+signed(MULTS_1_8(46)(PERCISION) & MULTS_1_8(46)(PERCISION downto 1));
			MULTS_2_4(47)<=signed(MULTS_1_7(47)(PERCISION) & MULTS_1_7(47)(PERCISION downto 1))+signed(MULTS_1_8(47)(PERCISION) & MULTS_1_8(47)(PERCISION downto 1));
			MULTS_2_4(48)<=signed(MULTS_1_7(48)(PERCISION) & MULTS_1_7(48)(PERCISION downto 1))+signed(MULTS_1_8(48)(PERCISION) & MULTS_1_8(48)(PERCISION downto 1));
			MULTS_2_4(49)<=signed(MULTS_1_7(49)(PERCISION) & MULTS_1_7(49)(PERCISION downto 1))+signed(MULTS_1_8(49)(PERCISION) & MULTS_1_8(49)(PERCISION downto 1));
			MULTS_2_4(50)<=signed(MULTS_1_7(50)(PERCISION) & MULTS_1_7(50)(PERCISION downto 1))+signed(MULTS_1_8(50)(PERCISION) & MULTS_1_8(50)(PERCISION downto 1));
			MULTS_2_4(51)<=signed(MULTS_1_7(51)(PERCISION) & MULTS_1_7(51)(PERCISION downto 1))+signed(MULTS_1_8(51)(PERCISION) & MULTS_1_8(51)(PERCISION downto 1));
			MULTS_2_4(52)<=signed(MULTS_1_7(52)(PERCISION) & MULTS_1_7(52)(PERCISION downto 1))+signed(MULTS_1_8(52)(PERCISION) & MULTS_1_8(52)(PERCISION downto 1));
			MULTS_2_4(53)<=signed(MULTS_1_7(53)(PERCISION) & MULTS_1_7(53)(PERCISION downto 1))+signed(MULTS_1_8(53)(PERCISION) & MULTS_1_8(53)(PERCISION downto 1));
			MULTS_2_4(54)<=signed(MULTS_1_7(54)(PERCISION) & MULTS_1_7(54)(PERCISION downto 1))+signed(MULTS_1_8(54)(PERCISION) & MULTS_1_8(54)(PERCISION downto 1));
			MULTS_2_4(55)<=signed(MULTS_1_7(55)(PERCISION) & MULTS_1_7(55)(PERCISION downto 1))+signed(MULTS_1_8(55)(PERCISION) & MULTS_1_8(55)(PERCISION downto 1));
			MULTS_2_4(56)<=signed(MULTS_1_7(56)(PERCISION) & MULTS_1_7(56)(PERCISION downto 1))+signed(MULTS_1_8(56)(PERCISION) & MULTS_1_8(56)(PERCISION downto 1));
			MULTS_2_4(57)<=signed(MULTS_1_7(57)(PERCISION) & MULTS_1_7(57)(PERCISION downto 1))+signed(MULTS_1_8(57)(PERCISION) & MULTS_1_8(57)(PERCISION downto 1));
			MULTS_2_4(58)<=signed(MULTS_1_7(58)(PERCISION) & MULTS_1_7(58)(PERCISION downto 1))+signed(MULTS_1_8(58)(PERCISION) & MULTS_1_8(58)(PERCISION downto 1));
			MULTS_2_4(59)<=signed(MULTS_1_7(59)(PERCISION) & MULTS_1_7(59)(PERCISION downto 1))+signed(MULTS_1_8(59)(PERCISION) & MULTS_1_8(59)(PERCISION downto 1));
			MULTS_2_4(60)<=signed(MULTS_1_7(60)(PERCISION) & MULTS_1_7(60)(PERCISION downto 1))+signed(MULTS_1_8(60)(PERCISION) & MULTS_1_8(60)(PERCISION downto 1));
			MULTS_2_4(61)<=signed(MULTS_1_7(61)(PERCISION) & MULTS_1_7(61)(PERCISION downto 1))+signed(MULTS_1_8(61)(PERCISION) & MULTS_1_8(61)(PERCISION downto 1));
			MULTS_2_4(62)<=signed(MULTS_1_7(62)(PERCISION) & MULTS_1_7(62)(PERCISION downto 1))+signed(MULTS_1_8(62)(PERCISION) & MULTS_1_8(62)(PERCISION downto 1));
			MULTS_2_4(63)<=signed(MULTS_1_7(63)(PERCISION) & MULTS_1_7(63)(PERCISION downto 1))+signed(MULTS_1_8(63)(PERCISION) & MULTS_1_8(63)(PERCISION downto 1));
			MULTS_2_4(64)<=signed(MULTS_1_7(64)(PERCISION) & MULTS_1_7(64)(PERCISION downto 1))+signed(MULTS_1_8(64)(PERCISION) & MULTS_1_8(64)(PERCISION downto 1));
			MULTS_2_4(65)<=signed(MULTS_1_7(65)(PERCISION) & MULTS_1_7(65)(PERCISION downto 1))+signed(MULTS_1_8(65)(PERCISION) & MULTS_1_8(65)(PERCISION downto 1));
			MULTS_2_4(66)<=signed(MULTS_1_7(66)(PERCISION) & MULTS_1_7(66)(PERCISION downto 1))+signed(MULTS_1_8(66)(PERCISION) & MULTS_1_8(66)(PERCISION downto 1));
			MULTS_2_4(67)<=signed(MULTS_1_7(67)(PERCISION) & MULTS_1_7(67)(PERCISION downto 1))+signed(MULTS_1_8(67)(PERCISION) & MULTS_1_8(67)(PERCISION downto 1));
			MULTS_2_4(68)<=signed(MULTS_1_7(68)(PERCISION) & MULTS_1_7(68)(PERCISION downto 1))+signed(MULTS_1_8(68)(PERCISION) & MULTS_1_8(68)(PERCISION downto 1));
			MULTS_2_4(69)<=signed(MULTS_1_7(69)(PERCISION) & MULTS_1_7(69)(PERCISION downto 1))+signed(MULTS_1_8(69)(PERCISION) & MULTS_1_8(69)(PERCISION downto 1));
			MULTS_2_4(70)<=signed(MULTS_1_7(70)(PERCISION) & MULTS_1_7(70)(PERCISION downto 1))+signed(MULTS_1_8(70)(PERCISION) & MULTS_1_8(70)(PERCISION downto 1));
			MULTS_2_4(71)<=signed(MULTS_1_7(71)(PERCISION) & MULTS_1_7(71)(PERCISION downto 1))+signed(MULTS_1_8(71)(PERCISION) & MULTS_1_8(71)(PERCISION downto 1));
			MULTS_2_4(72)<=signed(MULTS_1_7(72)(PERCISION) & MULTS_1_7(72)(PERCISION downto 1))+signed(MULTS_1_8(72)(PERCISION) & MULTS_1_8(72)(PERCISION downto 1));
			MULTS_2_4(73)<=signed(MULTS_1_7(73)(PERCISION) & MULTS_1_7(73)(PERCISION downto 1))+signed(MULTS_1_8(73)(PERCISION) & MULTS_1_8(73)(PERCISION downto 1));
			MULTS_2_4(74)<=signed(MULTS_1_7(74)(PERCISION) & MULTS_1_7(74)(PERCISION downto 1))+signed(MULTS_1_8(74)(PERCISION) & MULTS_1_8(74)(PERCISION downto 1));
			MULTS_2_4(75)<=signed(MULTS_1_7(75)(PERCISION) & MULTS_1_7(75)(PERCISION downto 1))+signed(MULTS_1_8(75)(PERCISION) & MULTS_1_8(75)(PERCISION downto 1));
			MULTS_2_4(76)<=signed(MULTS_1_7(76)(PERCISION) & MULTS_1_7(76)(PERCISION downto 1))+signed(MULTS_1_8(76)(PERCISION) & MULTS_1_8(76)(PERCISION downto 1));
			MULTS_2_4(77)<=signed(MULTS_1_7(77)(PERCISION) & MULTS_1_7(77)(PERCISION downto 1))+signed(MULTS_1_8(77)(PERCISION) & MULTS_1_8(77)(PERCISION downto 1));
			MULTS_2_4(78)<=signed(MULTS_1_7(78)(PERCISION) & MULTS_1_7(78)(PERCISION downto 1))+signed(MULTS_1_8(78)(PERCISION) & MULTS_1_8(78)(PERCISION downto 1));
			MULTS_2_4(79)<=signed(MULTS_1_7(79)(PERCISION) & MULTS_1_7(79)(PERCISION downto 1))+signed(MULTS_1_8(79)(PERCISION) & MULTS_1_8(79)(PERCISION downto 1));
			MULTS_2_4(80)<=signed(MULTS_1_7(80)(PERCISION) & MULTS_1_7(80)(PERCISION downto 1))+signed(MULTS_1_8(80)(PERCISION) & MULTS_1_8(80)(PERCISION downto 1));
			MULTS_2_4(81)<=signed(MULTS_1_7(81)(PERCISION) & MULTS_1_7(81)(PERCISION downto 1))+signed(MULTS_1_8(81)(PERCISION) & MULTS_1_8(81)(PERCISION downto 1));
			MULTS_2_4(82)<=signed(MULTS_1_7(82)(PERCISION) & MULTS_1_7(82)(PERCISION downto 1))+signed(MULTS_1_8(82)(PERCISION) & MULTS_1_8(82)(PERCISION downto 1));
			MULTS_2_4(83)<=signed(MULTS_1_7(83)(PERCISION) & MULTS_1_7(83)(PERCISION downto 1))+signed(MULTS_1_8(83)(PERCISION) & MULTS_1_8(83)(PERCISION downto 1));

			MULTS_2_5(0)<=signed(MULTS_1_9(0)(PERCISION) & MULTS_1_9(0)(PERCISION downto 1))+signed(MULTS_1_10(0)(PERCISION) & MULTS_1_10(0)(PERCISION downto 1));
			MULTS_2_5(1)<=signed(MULTS_1_9(1)(PERCISION) & MULTS_1_9(1)(PERCISION downto 1))+signed(MULTS_1_10(1)(PERCISION) & MULTS_1_10(1)(PERCISION downto 1));
			MULTS_2_5(2)<=signed(MULTS_1_9(2)(PERCISION) & MULTS_1_9(2)(PERCISION downto 1))+signed(MULTS_1_10(2)(PERCISION) & MULTS_1_10(2)(PERCISION downto 1));
			MULTS_2_5(3)<=signed(MULTS_1_9(3)(PERCISION) & MULTS_1_9(3)(PERCISION downto 1))+signed(MULTS_1_10(3)(PERCISION) & MULTS_1_10(3)(PERCISION downto 1));
			MULTS_2_5(4)<=signed(MULTS_1_9(4)(PERCISION) & MULTS_1_9(4)(PERCISION downto 1))+signed(MULTS_1_10(4)(PERCISION) & MULTS_1_10(4)(PERCISION downto 1));
			MULTS_2_5(5)<=signed(MULTS_1_9(5)(PERCISION) & MULTS_1_9(5)(PERCISION downto 1))+signed(MULTS_1_10(5)(PERCISION) & MULTS_1_10(5)(PERCISION downto 1));
			MULTS_2_5(6)<=signed(MULTS_1_9(6)(PERCISION) & MULTS_1_9(6)(PERCISION downto 1))+signed(MULTS_1_10(6)(PERCISION) & MULTS_1_10(6)(PERCISION downto 1));
			MULTS_2_5(7)<=signed(MULTS_1_9(7)(PERCISION) & MULTS_1_9(7)(PERCISION downto 1))+signed(MULTS_1_10(7)(PERCISION) & MULTS_1_10(7)(PERCISION downto 1));
			MULTS_2_5(8)<=signed(MULTS_1_9(8)(PERCISION) & MULTS_1_9(8)(PERCISION downto 1))+signed(MULTS_1_10(8)(PERCISION) & MULTS_1_10(8)(PERCISION downto 1));
			MULTS_2_5(9)<=signed(MULTS_1_9(9)(PERCISION) & MULTS_1_9(9)(PERCISION downto 1))+signed(MULTS_1_10(9)(PERCISION) & MULTS_1_10(9)(PERCISION downto 1));
			MULTS_2_5(10)<=signed(MULTS_1_9(10)(PERCISION) & MULTS_1_9(10)(PERCISION downto 1))+signed(MULTS_1_10(10)(PERCISION) & MULTS_1_10(10)(PERCISION downto 1));
			MULTS_2_5(11)<=signed(MULTS_1_9(11)(PERCISION) & MULTS_1_9(11)(PERCISION downto 1))+signed(MULTS_1_10(11)(PERCISION) & MULTS_1_10(11)(PERCISION downto 1));
			MULTS_2_5(12)<=signed(MULTS_1_9(12)(PERCISION) & MULTS_1_9(12)(PERCISION downto 1))+signed(MULTS_1_10(12)(PERCISION) & MULTS_1_10(12)(PERCISION downto 1));
			MULTS_2_5(13)<=signed(MULTS_1_9(13)(PERCISION) & MULTS_1_9(13)(PERCISION downto 1))+signed(MULTS_1_10(13)(PERCISION) & MULTS_1_10(13)(PERCISION downto 1));
			MULTS_2_5(14)<=signed(MULTS_1_9(14)(PERCISION) & MULTS_1_9(14)(PERCISION downto 1))+signed(MULTS_1_10(14)(PERCISION) & MULTS_1_10(14)(PERCISION downto 1));
			MULTS_2_5(15)<=signed(MULTS_1_9(15)(PERCISION) & MULTS_1_9(15)(PERCISION downto 1))+signed(MULTS_1_10(15)(PERCISION) & MULTS_1_10(15)(PERCISION downto 1));
			MULTS_2_5(16)<=signed(MULTS_1_9(16)(PERCISION) & MULTS_1_9(16)(PERCISION downto 1))+signed(MULTS_1_10(16)(PERCISION) & MULTS_1_10(16)(PERCISION downto 1));
			MULTS_2_5(17)<=signed(MULTS_1_9(17)(PERCISION) & MULTS_1_9(17)(PERCISION downto 1))+signed(MULTS_1_10(17)(PERCISION) & MULTS_1_10(17)(PERCISION downto 1));
			MULTS_2_5(18)<=signed(MULTS_1_9(18)(PERCISION) & MULTS_1_9(18)(PERCISION downto 1))+signed(MULTS_1_10(18)(PERCISION) & MULTS_1_10(18)(PERCISION downto 1));
			MULTS_2_5(19)<=signed(MULTS_1_9(19)(PERCISION) & MULTS_1_9(19)(PERCISION downto 1))+signed(MULTS_1_10(19)(PERCISION) & MULTS_1_10(19)(PERCISION downto 1));
			MULTS_2_5(20)<=signed(MULTS_1_9(20)(PERCISION) & MULTS_1_9(20)(PERCISION downto 1))+signed(MULTS_1_10(20)(PERCISION) & MULTS_1_10(20)(PERCISION downto 1));
			MULTS_2_5(21)<=signed(MULTS_1_9(21)(PERCISION) & MULTS_1_9(21)(PERCISION downto 1))+signed(MULTS_1_10(21)(PERCISION) & MULTS_1_10(21)(PERCISION downto 1));
			MULTS_2_5(22)<=signed(MULTS_1_9(22)(PERCISION) & MULTS_1_9(22)(PERCISION downto 1))+signed(MULTS_1_10(22)(PERCISION) & MULTS_1_10(22)(PERCISION downto 1));
			MULTS_2_5(23)<=signed(MULTS_1_9(23)(PERCISION) & MULTS_1_9(23)(PERCISION downto 1))+signed(MULTS_1_10(23)(PERCISION) & MULTS_1_10(23)(PERCISION downto 1));
			MULTS_2_5(24)<=signed(MULTS_1_9(24)(PERCISION) & MULTS_1_9(24)(PERCISION downto 1))+signed(MULTS_1_10(24)(PERCISION) & MULTS_1_10(24)(PERCISION downto 1));
			MULTS_2_5(25)<=signed(MULTS_1_9(25)(PERCISION) & MULTS_1_9(25)(PERCISION downto 1))+signed(MULTS_1_10(25)(PERCISION) & MULTS_1_10(25)(PERCISION downto 1));
			MULTS_2_5(26)<=signed(MULTS_1_9(26)(PERCISION) & MULTS_1_9(26)(PERCISION downto 1))+signed(MULTS_1_10(26)(PERCISION) & MULTS_1_10(26)(PERCISION downto 1));
			MULTS_2_5(27)<=signed(MULTS_1_9(27)(PERCISION) & MULTS_1_9(27)(PERCISION downto 1))+signed(MULTS_1_10(27)(PERCISION) & MULTS_1_10(27)(PERCISION downto 1));
			MULTS_2_5(28)<=signed(MULTS_1_9(28)(PERCISION) & MULTS_1_9(28)(PERCISION downto 1))+signed(MULTS_1_10(28)(PERCISION) & MULTS_1_10(28)(PERCISION downto 1));
			MULTS_2_5(29)<=signed(MULTS_1_9(29)(PERCISION) & MULTS_1_9(29)(PERCISION downto 1))+signed(MULTS_1_10(29)(PERCISION) & MULTS_1_10(29)(PERCISION downto 1));
			MULTS_2_5(30)<=signed(MULTS_1_9(30)(PERCISION) & MULTS_1_9(30)(PERCISION downto 1))+signed(MULTS_1_10(30)(PERCISION) & MULTS_1_10(30)(PERCISION downto 1));
			MULTS_2_5(31)<=signed(MULTS_1_9(31)(PERCISION) & MULTS_1_9(31)(PERCISION downto 1))+signed(MULTS_1_10(31)(PERCISION) & MULTS_1_10(31)(PERCISION downto 1));
			MULTS_2_5(32)<=signed(MULTS_1_9(32)(PERCISION) & MULTS_1_9(32)(PERCISION downto 1))+signed(MULTS_1_10(32)(PERCISION) & MULTS_1_10(32)(PERCISION downto 1));
			MULTS_2_5(33)<=signed(MULTS_1_9(33)(PERCISION) & MULTS_1_9(33)(PERCISION downto 1))+signed(MULTS_1_10(33)(PERCISION) & MULTS_1_10(33)(PERCISION downto 1));
			MULTS_2_5(34)<=signed(MULTS_1_9(34)(PERCISION) & MULTS_1_9(34)(PERCISION downto 1))+signed(MULTS_1_10(34)(PERCISION) & MULTS_1_10(34)(PERCISION downto 1));
			MULTS_2_5(35)<=signed(MULTS_1_9(35)(PERCISION) & MULTS_1_9(35)(PERCISION downto 1))+signed(MULTS_1_10(35)(PERCISION) & MULTS_1_10(35)(PERCISION downto 1));
			MULTS_2_5(36)<=signed(MULTS_1_9(36)(PERCISION) & MULTS_1_9(36)(PERCISION downto 1))+signed(MULTS_1_10(36)(PERCISION) & MULTS_1_10(36)(PERCISION downto 1));
			MULTS_2_5(37)<=signed(MULTS_1_9(37)(PERCISION) & MULTS_1_9(37)(PERCISION downto 1))+signed(MULTS_1_10(37)(PERCISION) & MULTS_1_10(37)(PERCISION downto 1));
			MULTS_2_5(38)<=signed(MULTS_1_9(38)(PERCISION) & MULTS_1_9(38)(PERCISION downto 1))+signed(MULTS_1_10(38)(PERCISION) & MULTS_1_10(38)(PERCISION downto 1));
			MULTS_2_5(39)<=signed(MULTS_1_9(39)(PERCISION) & MULTS_1_9(39)(PERCISION downto 1))+signed(MULTS_1_10(39)(PERCISION) & MULTS_1_10(39)(PERCISION downto 1));
			MULTS_2_5(40)<=signed(MULTS_1_9(40)(PERCISION) & MULTS_1_9(40)(PERCISION downto 1))+signed(MULTS_1_10(40)(PERCISION) & MULTS_1_10(40)(PERCISION downto 1));
			MULTS_2_5(41)<=signed(MULTS_1_9(41)(PERCISION) & MULTS_1_9(41)(PERCISION downto 1))+signed(MULTS_1_10(41)(PERCISION) & MULTS_1_10(41)(PERCISION downto 1));
			MULTS_2_5(42)<=signed(MULTS_1_9(42)(PERCISION) & MULTS_1_9(42)(PERCISION downto 1))+signed(MULTS_1_10(42)(PERCISION) & MULTS_1_10(42)(PERCISION downto 1));
			MULTS_2_5(43)<=signed(MULTS_1_9(43)(PERCISION) & MULTS_1_9(43)(PERCISION downto 1))+signed(MULTS_1_10(43)(PERCISION) & MULTS_1_10(43)(PERCISION downto 1));
			MULTS_2_5(44)<=signed(MULTS_1_9(44)(PERCISION) & MULTS_1_9(44)(PERCISION downto 1))+signed(MULTS_1_10(44)(PERCISION) & MULTS_1_10(44)(PERCISION downto 1));
			MULTS_2_5(45)<=signed(MULTS_1_9(45)(PERCISION) & MULTS_1_9(45)(PERCISION downto 1))+signed(MULTS_1_10(45)(PERCISION) & MULTS_1_10(45)(PERCISION downto 1));
			MULTS_2_5(46)<=signed(MULTS_1_9(46)(PERCISION) & MULTS_1_9(46)(PERCISION downto 1))+signed(MULTS_1_10(46)(PERCISION) & MULTS_1_10(46)(PERCISION downto 1));
			MULTS_2_5(47)<=signed(MULTS_1_9(47)(PERCISION) & MULTS_1_9(47)(PERCISION downto 1))+signed(MULTS_1_10(47)(PERCISION) & MULTS_1_10(47)(PERCISION downto 1));
			MULTS_2_5(48)<=signed(MULTS_1_9(48)(PERCISION) & MULTS_1_9(48)(PERCISION downto 1))+signed(MULTS_1_10(48)(PERCISION) & MULTS_1_10(48)(PERCISION downto 1));
			MULTS_2_5(49)<=signed(MULTS_1_9(49)(PERCISION) & MULTS_1_9(49)(PERCISION downto 1))+signed(MULTS_1_10(49)(PERCISION) & MULTS_1_10(49)(PERCISION downto 1));
			MULTS_2_5(50)<=signed(MULTS_1_9(50)(PERCISION) & MULTS_1_9(50)(PERCISION downto 1))+signed(MULTS_1_10(50)(PERCISION) & MULTS_1_10(50)(PERCISION downto 1));
			MULTS_2_5(51)<=signed(MULTS_1_9(51)(PERCISION) & MULTS_1_9(51)(PERCISION downto 1))+signed(MULTS_1_10(51)(PERCISION) & MULTS_1_10(51)(PERCISION downto 1));
			MULTS_2_5(52)<=signed(MULTS_1_9(52)(PERCISION) & MULTS_1_9(52)(PERCISION downto 1))+signed(MULTS_1_10(52)(PERCISION) & MULTS_1_10(52)(PERCISION downto 1));
			MULTS_2_5(53)<=signed(MULTS_1_9(53)(PERCISION) & MULTS_1_9(53)(PERCISION downto 1))+signed(MULTS_1_10(53)(PERCISION) & MULTS_1_10(53)(PERCISION downto 1));
			MULTS_2_5(54)<=signed(MULTS_1_9(54)(PERCISION) & MULTS_1_9(54)(PERCISION downto 1))+signed(MULTS_1_10(54)(PERCISION) & MULTS_1_10(54)(PERCISION downto 1));
			MULTS_2_5(55)<=signed(MULTS_1_9(55)(PERCISION) & MULTS_1_9(55)(PERCISION downto 1))+signed(MULTS_1_10(55)(PERCISION) & MULTS_1_10(55)(PERCISION downto 1));
			MULTS_2_5(56)<=signed(MULTS_1_9(56)(PERCISION) & MULTS_1_9(56)(PERCISION downto 1))+signed(MULTS_1_10(56)(PERCISION) & MULTS_1_10(56)(PERCISION downto 1));
			MULTS_2_5(57)<=signed(MULTS_1_9(57)(PERCISION) & MULTS_1_9(57)(PERCISION downto 1))+signed(MULTS_1_10(57)(PERCISION) & MULTS_1_10(57)(PERCISION downto 1));
			MULTS_2_5(58)<=signed(MULTS_1_9(58)(PERCISION) & MULTS_1_9(58)(PERCISION downto 1))+signed(MULTS_1_10(58)(PERCISION) & MULTS_1_10(58)(PERCISION downto 1));
			MULTS_2_5(59)<=signed(MULTS_1_9(59)(PERCISION) & MULTS_1_9(59)(PERCISION downto 1))+signed(MULTS_1_10(59)(PERCISION) & MULTS_1_10(59)(PERCISION downto 1));
			MULTS_2_5(60)<=signed(MULTS_1_9(60)(PERCISION) & MULTS_1_9(60)(PERCISION downto 1))+signed(MULTS_1_10(60)(PERCISION) & MULTS_1_10(60)(PERCISION downto 1));
			MULTS_2_5(61)<=signed(MULTS_1_9(61)(PERCISION) & MULTS_1_9(61)(PERCISION downto 1))+signed(MULTS_1_10(61)(PERCISION) & MULTS_1_10(61)(PERCISION downto 1));
			MULTS_2_5(62)<=signed(MULTS_1_9(62)(PERCISION) & MULTS_1_9(62)(PERCISION downto 1))+signed(MULTS_1_10(62)(PERCISION) & MULTS_1_10(62)(PERCISION downto 1));
			MULTS_2_5(63)<=signed(MULTS_1_9(63)(PERCISION) & MULTS_1_9(63)(PERCISION downto 1))+signed(MULTS_1_10(63)(PERCISION) & MULTS_1_10(63)(PERCISION downto 1));
			MULTS_2_5(64)<=signed(MULTS_1_9(64)(PERCISION) & MULTS_1_9(64)(PERCISION downto 1))+signed(MULTS_1_10(64)(PERCISION) & MULTS_1_10(64)(PERCISION downto 1));
			MULTS_2_5(65)<=signed(MULTS_1_9(65)(PERCISION) & MULTS_1_9(65)(PERCISION downto 1))+signed(MULTS_1_10(65)(PERCISION) & MULTS_1_10(65)(PERCISION downto 1));
			MULTS_2_5(66)<=signed(MULTS_1_9(66)(PERCISION) & MULTS_1_9(66)(PERCISION downto 1))+signed(MULTS_1_10(66)(PERCISION) & MULTS_1_10(66)(PERCISION downto 1));
			MULTS_2_5(67)<=signed(MULTS_1_9(67)(PERCISION) & MULTS_1_9(67)(PERCISION downto 1))+signed(MULTS_1_10(67)(PERCISION) & MULTS_1_10(67)(PERCISION downto 1));
			MULTS_2_5(68)<=signed(MULTS_1_9(68)(PERCISION) & MULTS_1_9(68)(PERCISION downto 1))+signed(MULTS_1_10(68)(PERCISION) & MULTS_1_10(68)(PERCISION downto 1));
			MULTS_2_5(69)<=signed(MULTS_1_9(69)(PERCISION) & MULTS_1_9(69)(PERCISION downto 1))+signed(MULTS_1_10(69)(PERCISION) & MULTS_1_10(69)(PERCISION downto 1));
			MULTS_2_5(70)<=signed(MULTS_1_9(70)(PERCISION) & MULTS_1_9(70)(PERCISION downto 1))+signed(MULTS_1_10(70)(PERCISION) & MULTS_1_10(70)(PERCISION downto 1));
			MULTS_2_5(71)<=signed(MULTS_1_9(71)(PERCISION) & MULTS_1_9(71)(PERCISION downto 1))+signed(MULTS_1_10(71)(PERCISION) & MULTS_1_10(71)(PERCISION downto 1));
			MULTS_2_5(72)<=signed(MULTS_1_9(72)(PERCISION) & MULTS_1_9(72)(PERCISION downto 1))+signed(MULTS_1_10(72)(PERCISION) & MULTS_1_10(72)(PERCISION downto 1));
			MULTS_2_5(73)<=signed(MULTS_1_9(73)(PERCISION) & MULTS_1_9(73)(PERCISION downto 1))+signed(MULTS_1_10(73)(PERCISION) & MULTS_1_10(73)(PERCISION downto 1));
			MULTS_2_5(74)<=signed(MULTS_1_9(74)(PERCISION) & MULTS_1_9(74)(PERCISION downto 1))+signed(MULTS_1_10(74)(PERCISION) & MULTS_1_10(74)(PERCISION downto 1));
			MULTS_2_5(75)<=signed(MULTS_1_9(75)(PERCISION) & MULTS_1_9(75)(PERCISION downto 1))+signed(MULTS_1_10(75)(PERCISION) & MULTS_1_10(75)(PERCISION downto 1));
			MULTS_2_5(76)<=signed(MULTS_1_9(76)(PERCISION) & MULTS_1_9(76)(PERCISION downto 1))+signed(MULTS_1_10(76)(PERCISION) & MULTS_1_10(76)(PERCISION downto 1));
			MULTS_2_5(77)<=signed(MULTS_1_9(77)(PERCISION) & MULTS_1_9(77)(PERCISION downto 1))+signed(MULTS_1_10(77)(PERCISION) & MULTS_1_10(77)(PERCISION downto 1));
			MULTS_2_5(78)<=signed(MULTS_1_9(78)(PERCISION) & MULTS_1_9(78)(PERCISION downto 1))+signed(MULTS_1_10(78)(PERCISION) & MULTS_1_10(78)(PERCISION downto 1));
			MULTS_2_5(79)<=signed(MULTS_1_9(79)(PERCISION) & MULTS_1_9(79)(PERCISION downto 1))+signed(MULTS_1_10(79)(PERCISION) & MULTS_1_10(79)(PERCISION downto 1));
			MULTS_2_5(80)<=signed(MULTS_1_9(80)(PERCISION) & MULTS_1_9(80)(PERCISION downto 1))+signed(MULTS_1_10(80)(PERCISION) & MULTS_1_10(80)(PERCISION downto 1));
			MULTS_2_5(81)<=signed(MULTS_1_9(81)(PERCISION) & MULTS_1_9(81)(PERCISION downto 1))+signed(MULTS_1_10(81)(PERCISION) & MULTS_1_10(81)(PERCISION downto 1));
			MULTS_2_5(82)<=signed(MULTS_1_9(82)(PERCISION) & MULTS_1_9(82)(PERCISION downto 1))+signed(MULTS_1_10(82)(PERCISION) & MULTS_1_10(82)(PERCISION downto 1));
			MULTS_2_5(83)<=signed(MULTS_1_9(83)(PERCISION) & MULTS_1_9(83)(PERCISION downto 1))+signed(MULTS_1_10(83)(PERCISION) & MULTS_1_10(83)(PERCISION downto 1));

			MULTS_2_6(0)<=signed(MULTS_1_11(0)(PERCISION) & MULTS_1_11(0)(PERCISION downto 1))+signed(MULTS_1_12(0)(PERCISION) & MULTS_1_12(0)(PERCISION downto 1));
			MULTS_2_6(1)<=signed(MULTS_1_11(1)(PERCISION) & MULTS_1_11(1)(PERCISION downto 1))+signed(MULTS_1_12(1)(PERCISION) & MULTS_1_12(1)(PERCISION downto 1));
			MULTS_2_6(2)<=signed(MULTS_1_11(2)(PERCISION) & MULTS_1_11(2)(PERCISION downto 1))+signed(MULTS_1_12(2)(PERCISION) & MULTS_1_12(2)(PERCISION downto 1));
			MULTS_2_6(3)<=signed(MULTS_1_11(3)(PERCISION) & MULTS_1_11(3)(PERCISION downto 1))+signed(MULTS_1_12(3)(PERCISION) & MULTS_1_12(3)(PERCISION downto 1));
			MULTS_2_6(4)<=signed(MULTS_1_11(4)(PERCISION) & MULTS_1_11(4)(PERCISION downto 1))+signed(MULTS_1_12(4)(PERCISION) & MULTS_1_12(4)(PERCISION downto 1));
			MULTS_2_6(5)<=signed(MULTS_1_11(5)(PERCISION) & MULTS_1_11(5)(PERCISION downto 1))+signed(MULTS_1_12(5)(PERCISION) & MULTS_1_12(5)(PERCISION downto 1));
			MULTS_2_6(6)<=signed(MULTS_1_11(6)(PERCISION) & MULTS_1_11(6)(PERCISION downto 1))+signed(MULTS_1_12(6)(PERCISION) & MULTS_1_12(6)(PERCISION downto 1));
			MULTS_2_6(7)<=signed(MULTS_1_11(7)(PERCISION) & MULTS_1_11(7)(PERCISION downto 1))+signed(MULTS_1_12(7)(PERCISION) & MULTS_1_12(7)(PERCISION downto 1));
			MULTS_2_6(8)<=signed(MULTS_1_11(8)(PERCISION) & MULTS_1_11(8)(PERCISION downto 1))+signed(MULTS_1_12(8)(PERCISION) & MULTS_1_12(8)(PERCISION downto 1));
			MULTS_2_6(9)<=signed(MULTS_1_11(9)(PERCISION) & MULTS_1_11(9)(PERCISION downto 1))+signed(MULTS_1_12(9)(PERCISION) & MULTS_1_12(9)(PERCISION downto 1));
			MULTS_2_6(10)<=signed(MULTS_1_11(10)(PERCISION) & MULTS_1_11(10)(PERCISION downto 1))+signed(MULTS_1_12(10)(PERCISION) & MULTS_1_12(10)(PERCISION downto 1));
			MULTS_2_6(11)<=signed(MULTS_1_11(11)(PERCISION) & MULTS_1_11(11)(PERCISION downto 1))+signed(MULTS_1_12(11)(PERCISION) & MULTS_1_12(11)(PERCISION downto 1));
			MULTS_2_6(12)<=signed(MULTS_1_11(12)(PERCISION) & MULTS_1_11(12)(PERCISION downto 1))+signed(MULTS_1_12(12)(PERCISION) & MULTS_1_12(12)(PERCISION downto 1));
			MULTS_2_6(13)<=signed(MULTS_1_11(13)(PERCISION) & MULTS_1_11(13)(PERCISION downto 1))+signed(MULTS_1_12(13)(PERCISION) & MULTS_1_12(13)(PERCISION downto 1));
			MULTS_2_6(14)<=signed(MULTS_1_11(14)(PERCISION) & MULTS_1_11(14)(PERCISION downto 1))+signed(MULTS_1_12(14)(PERCISION) & MULTS_1_12(14)(PERCISION downto 1));
			MULTS_2_6(15)<=signed(MULTS_1_11(15)(PERCISION) & MULTS_1_11(15)(PERCISION downto 1))+signed(MULTS_1_12(15)(PERCISION) & MULTS_1_12(15)(PERCISION downto 1));
			MULTS_2_6(16)<=signed(MULTS_1_11(16)(PERCISION) & MULTS_1_11(16)(PERCISION downto 1))+signed(MULTS_1_12(16)(PERCISION) & MULTS_1_12(16)(PERCISION downto 1));
			MULTS_2_6(17)<=signed(MULTS_1_11(17)(PERCISION) & MULTS_1_11(17)(PERCISION downto 1))+signed(MULTS_1_12(17)(PERCISION) & MULTS_1_12(17)(PERCISION downto 1));
			MULTS_2_6(18)<=signed(MULTS_1_11(18)(PERCISION) & MULTS_1_11(18)(PERCISION downto 1))+signed(MULTS_1_12(18)(PERCISION) & MULTS_1_12(18)(PERCISION downto 1));
			MULTS_2_6(19)<=signed(MULTS_1_11(19)(PERCISION) & MULTS_1_11(19)(PERCISION downto 1))+signed(MULTS_1_12(19)(PERCISION) & MULTS_1_12(19)(PERCISION downto 1));
			MULTS_2_6(20)<=signed(MULTS_1_11(20)(PERCISION) & MULTS_1_11(20)(PERCISION downto 1))+signed(MULTS_1_12(20)(PERCISION) & MULTS_1_12(20)(PERCISION downto 1));
			MULTS_2_6(21)<=signed(MULTS_1_11(21)(PERCISION) & MULTS_1_11(21)(PERCISION downto 1))+signed(MULTS_1_12(21)(PERCISION) & MULTS_1_12(21)(PERCISION downto 1));
			MULTS_2_6(22)<=signed(MULTS_1_11(22)(PERCISION) & MULTS_1_11(22)(PERCISION downto 1))+signed(MULTS_1_12(22)(PERCISION) & MULTS_1_12(22)(PERCISION downto 1));
			MULTS_2_6(23)<=signed(MULTS_1_11(23)(PERCISION) & MULTS_1_11(23)(PERCISION downto 1))+signed(MULTS_1_12(23)(PERCISION) & MULTS_1_12(23)(PERCISION downto 1));
			MULTS_2_6(24)<=signed(MULTS_1_11(24)(PERCISION) & MULTS_1_11(24)(PERCISION downto 1))+signed(MULTS_1_12(24)(PERCISION) & MULTS_1_12(24)(PERCISION downto 1));
			MULTS_2_6(25)<=signed(MULTS_1_11(25)(PERCISION) & MULTS_1_11(25)(PERCISION downto 1))+signed(MULTS_1_12(25)(PERCISION) & MULTS_1_12(25)(PERCISION downto 1));
			MULTS_2_6(26)<=signed(MULTS_1_11(26)(PERCISION) & MULTS_1_11(26)(PERCISION downto 1))+signed(MULTS_1_12(26)(PERCISION) & MULTS_1_12(26)(PERCISION downto 1));
			MULTS_2_6(27)<=signed(MULTS_1_11(27)(PERCISION) & MULTS_1_11(27)(PERCISION downto 1))+signed(MULTS_1_12(27)(PERCISION) & MULTS_1_12(27)(PERCISION downto 1));
			MULTS_2_6(28)<=signed(MULTS_1_11(28)(PERCISION) & MULTS_1_11(28)(PERCISION downto 1))+signed(MULTS_1_12(28)(PERCISION) & MULTS_1_12(28)(PERCISION downto 1));
			MULTS_2_6(29)<=signed(MULTS_1_11(29)(PERCISION) & MULTS_1_11(29)(PERCISION downto 1))+signed(MULTS_1_12(29)(PERCISION) & MULTS_1_12(29)(PERCISION downto 1));
			MULTS_2_6(30)<=signed(MULTS_1_11(30)(PERCISION) & MULTS_1_11(30)(PERCISION downto 1))+signed(MULTS_1_12(30)(PERCISION) & MULTS_1_12(30)(PERCISION downto 1));
			MULTS_2_6(31)<=signed(MULTS_1_11(31)(PERCISION) & MULTS_1_11(31)(PERCISION downto 1))+signed(MULTS_1_12(31)(PERCISION) & MULTS_1_12(31)(PERCISION downto 1));
			MULTS_2_6(32)<=signed(MULTS_1_11(32)(PERCISION) & MULTS_1_11(32)(PERCISION downto 1))+signed(MULTS_1_12(32)(PERCISION) & MULTS_1_12(32)(PERCISION downto 1));
			MULTS_2_6(33)<=signed(MULTS_1_11(33)(PERCISION) & MULTS_1_11(33)(PERCISION downto 1))+signed(MULTS_1_12(33)(PERCISION) & MULTS_1_12(33)(PERCISION downto 1));
			MULTS_2_6(34)<=signed(MULTS_1_11(34)(PERCISION) & MULTS_1_11(34)(PERCISION downto 1))+signed(MULTS_1_12(34)(PERCISION) & MULTS_1_12(34)(PERCISION downto 1));
			MULTS_2_6(35)<=signed(MULTS_1_11(35)(PERCISION) & MULTS_1_11(35)(PERCISION downto 1))+signed(MULTS_1_12(35)(PERCISION) & MULTS_1_12(35)(PERCISION downto 1));
			MULTS_2_6(36)<=signed(MULTS_1_11(36)(PERCISION) & MULTS_1_11(36)(PERCISION downto 1))+signed(MULTS_1_12(36)(PERCISION) & MULTS_1_12(36)(PERCISION downto 1));
			MULTS_2_6(37)<=signed(MULTS_1_11(37)(PERCISION) & MULTS_1_11(37)(PERCISION downto 1))+signed(MULTS_1_12(37)(PERCISION) & MULTS_1_12(37)(PERCISION downto 1));
			MULTS_2_6(38)<=signed(MULTS_1_11(38)(PERCISION) & MULTS_1_11(38)(PERCISION downto 1))+signed(MULTS_1_12(38)(PERCISION) & MULTS_1_12(38)(PERCISION downto 1));
			MULTS_2_6(39)<=signed(MULTS_1_11(39)(PERCISION) & MULTS_1_11(39)(PERCISION downto 1))+signed(MULTS_1_12(39)(PERCISION) & MULTS_1_12(39)(PERCISION downto 1));
			MULTS_2_6(40)<=signed(MULTS_1_11(40)(PERCISION) & MULTS_1_11(40)(PERCISION downto 1))+signed(MULTS_1_12(40)(PERCISION) & MULTS_1_12(40)(PERCISION downto 1));
			MULTS_2_6(41)<=signed(MULTS_1_11(41)(PERCISION) & MULTS_1_11(41)(PERCISION downto 1))+signed(MULTS_1_12(41)(PERCISION) & MULTS_1_12(41)(PERCISION downto 1));
			MULTS_2_6(42)<=signed(MULTS_1_11(42)(PERCISION) & MULTS_1_11(42)(PERCISION downto 1))+signed(MULTS_1_12(42)(PERCISION) & MULTS_1_12(42)(PERCISION downto 1));
			MULTS_2_6(43)<=signed(MULTS_1_11(43)(PERCISION) & MULTS_1_11(43)(PERCISION downto 1))+signed(MULTS_1_12(43)(PERCISION) & MULTS_1_12(43)(PERCISION downto 1));
			MULTS_2_6(44)<=signed(MULTS_1_11(44)(PERCISION) & MULTS_1_11(44)(PERCISION downto 1))+signed(MULTS_1_12(44)(PERCISION) & MULTS_1_12(44)(PERCISION downto 1));
			MULTS_2_6(45)<=signed(MULTS_1_11(45)(PERCISION) & MULTS_1_11(45)(PERCISION downto 1))+signed(MULTS_1_12(45)(PERCISION) & MULTS_1_12(45)(PERCISION downto 1));
			MULTS_2_6(46)<=signed(MULTS_1_11(46)(PERCISION) & MULTS_1_11(46)(PERCISION downto 1))+signed(MULTS_1_12(46)(PERCISION) & MULTS_1_12(46)(PERCISION downto 1));
			MULTS_2_6(47)<=signed(MULTS_1_11(47)(PERCISION) & MULTS_1_11(47)(PERCISION downto 1))+signed(MULTS_1_12(47)(PERCISION) & MULTS_1_12(47)(PERCISION downto 1));
			MULTS_2_6(48)<=signed(MULTS_1_11(48)(PERCISION) & MULTS_1_11(48)(PERCISION downto 1))+signed(MULTS_1_12(48)(PERCISION) & MULTS_1_12(48)(PERCISION downto 1));
			MULTS_2_6(49)<=signed(MULTS_1_11(49)(PERCISION) & MULTS_1_11(49)(PERCISION downto 1))+signed(MULTS_1_12(49)(PERCISION) & MULTS_1_12(49)(PERCISION downto 1));
			MULTS_2_6(50)<=signed(MULTS_1_11(50)(PERCISION) & MULTS_1_11(50)(PERCISION downto 1))+signed(MULTS_1_12(50)(PERCISION) & MULTS_1_12(50)(PERCISION downto 1));
			MULTS_2_6(51)<=signed(MULTS_1_11(51)(PERCISION) & MULTS_1_11(51)(PERCISION downto 1))+signed(MULTS_1_12(51)(PERCISION) & MULTS_1_12(51)(PERCISION downto 1));
			MULTS_2_6(52)<=signed(MULTS_1_11(52)(PERCISION) & MULTS_1_11(52)(PERCISION downto 1))+signed(MULTS_1_12(52)(PERCISION) & MULTS_1_12(52)(PERCISION downto 1));
			MULTS_2_6(53)<=signed(MULTS_1_11(53)(PERCISION) & MULTS_1_11(53)(PERCISION downto 1))+signed(MULTS_1_12(53)(PERCISION) & MULTS_1_12(53)(PERCISION downto 1));
			MULTS_2_6(54)<=signed(MULTS_1_11(54)(PERCISION) & MULTS_1_11(54)(PERCISION downto 1))+signed(MULTS_1_12(54)(PERCISION) & MULTS_1_12(54)(PERCISION downto 1));
			MULTS_2_6(55)<=signed(MULTS_1_11(55)(PERCISION) & MULTS_1_11(55)(PERCISION downto 1))+signed(MULTS_1_12(55)(PERCISION) & MULTS_1_12(55)(PERCISION downto 1));
			MULTS_2_6(56)<=signed(MULTS_1_11(56)(PERCISION) & MULTS_1_11(56)(PERCISION downto 1))+signed(MULTS_1_12(56)(PERCISION) & MULTS_1_12(56)(PERCISION downto 1));
			MULTS_2_6(57)<=signed(MULTS_1_11(57)(PERCISION) & MULTS_1_11(57)(PERCISION downto 1))+signed(MULTS_1_12(57)(PERCISION) & MULTS_1_12(57)(PERCISION downto 1));
			MULTS_2_6(58)<=signed(MULTS_1_11(58)(PERCISION) & MULTS_1_11(58)(PERCISION downto 1))+signed(MULTS_1_12(58)(PERCISION) & MULTS_1_12(58)(PERCISION downto 1));
			MULTS_2_6(59)<=signed(MULTS_1_11(59)(PERCISION) & MULTS_1_11(59)(PERCISION downto 1))+signed(MULTS_1_12(59)(PERCISION) & MULTS_1_12(59)(PERCISION downto 1));
			MULTS_2_6(60)<=signed(MULTS_1_11(60)(PERCISION) & MULTS_1_11(60)(PERCISION downto 1))+signed(MULTS_1_12(60)(PERCISION) & MULTS_1_12(60)(PERCISION downto 1));
			MULTS_2_6(61)<=signed(MULTS_1_11(61)(PERCISION) & MULTS_1_11(61)(PERCISION downto 1))+signed(MULTS_1_12(61)(PERCISION) & MULTS_1_12(61)(PERCISION downto 1));
			MULTS_2_6(62)<=signed(MULTS_1_11(62)(PERCISION) & MULTS_1_11(62)(PERCISION downto 1))+signed(MULTS_1_12(62)(PERCISION) & MULTS_1_12(62)(PERCISION downto 1));
			MULTS_2_6(63)<=signed(MULTS_1_11(63)(PERCISION) & MULTS_1_11(63)(PERCISION downto 1))+signed(MULTS_1_12(63)(PERCISION) & MULTS_1_12(63)(PERCISION downto 1));
			MULTS_2_6(64)<=signed(MULTS_1_11(64)(PERCISION) & MULTS_1_11(64)(PERCISION downto 1))+signed(MULTS_1_12(64)(PERCISION) & MULTS_1_12(64)(PERCISION downto 1));
			MULTS_2_6(65)<=signed(MULTS_1_11(65)(PERCISION) & MULTS_1_11(65)(PERCISION downto 1))+signed(MULTS_1_12(65)(PERCISION) & MULTS_1_12(65)(PERCISION downto 1));
			MULTS_2_6(66)<=signed(MULTS_1_11(66)(PERCISION) & MULTS_1_11(66)(PERCISION downto 1))+signed(MULTS_1_12(66)(PERCISION) & MULTS_1_12(66)(PERCISION downto 1));
			MULTS_2_6(67)<=signed(MULTS_1_11(67)(PERCISION) & MULTS_1_11(67)(PERCISION downto 1))+signed(MULTS_1_12(67)(PERCISION) & MULTS_1_12(67)(PERCISION downto 1));
			MULTS_2_6(68)<=signed(MULTS_1_11(68)(PERCISION) & MULTS_1_11(68)(PERCISION downto 1))+signed(MULTS_1_12(68)(PERCISION) & MULTS_1_12(68)(PERCISION downto 1));
			MULTS_2_6(69)<=signed(MULTS_1_11(69)(PERCISION) & MULTS_1_11(69)(PERCISION downto 1))+signed(MULTS_1_12(69)(PERCISION) & MULTS_1_12(69)(PERCISION downto 1));
			MULTS_2_6(70)<=signed(MULTS_1_11(70)(PERCISION) & MULTS_1_11(70)(PERCISION downto 1))+signed(MULTS_1_12(70)(PERCISION) & MULTS_1_12(70)(PERCISION downto 1));
			MULTS_2_6(71)<=signed(MULTS_1_11(71)(PERCISION) & MULTS_1_11(71)(PERCISION downto 1))+signed(MULTS_1_12(71)(PERCISION) & MULTS_1_12(71)(PERCISION downto 1));
			MULTS_2_6(72)<=signed(MULTS_1_11(72)(PERCISION) & MULTS_1_11(72)(PERCISION downto 1))+signed(MULTS_1_12(72)(PERCISION) & MULTS_1_12(72)(PERCISION downto 1));
			MULTS_2_6(73)<=signed(MULTS_1_11(73)(PERCISION) & MULTS_1_11(73)(PERCISION downto 1))+signed(MULTS_1_12(73)(PERCISION) & MULTS_1_12(73)(PERCISION downto 1));
			MULTS_2_6(74)<=signed(MULTS_1_11(74)(PERCISION) & MULTS_1_11(74)(PERCISION downto 1))+signed(MULTS_1_12(74)(PERCISION) & MULTS_1_12(74)(PERCISION downto 1));
			MULTS_2_6(75)<=signed(MULTS_1_11(75)(PERCISION) & MULTS_1_11(75)(PERCISION downto 1))+signed(MULTS_1_12(75)(PERCISION) & MULTS_1_12(75)(PERCISION downto 1));
			MULTS_2_6(76)<=signed(MULTS_1_11(76)(PERCISION) & MULTS_1_11(76)(PERCISION downto 1))+signed(MULTS_1_12(76)(PERCISION) & MULTS_1_12(76)(PERCISION downto 1));
			MULTS_2_6(77)<=signed(MULTS_1_11(77)(PERCISION) & MULTS_1_11(77)(PERCISION downto 1))+signed(MULTS_1_12(77)(PERCISION) & MULTS_1_12(77)(PERCISION downto 1));
			MULTS_2_6(78)<=signed(MULTS_1_11(78)(PERCISION) & MULTS_1_11(78)(PERCISION downto 1))+signed(MULTS_1_12(78)(PERCISION) & MULTS_1_12(78)(PERCISION downto 1));
			MULTS_2_6(79)<=signed(MULTS_1_11(79)(PERCISION) & MULTS_1_11(79)(PERCISION downto 1))+signed(MULTS_1_12(79)(PERCISION) & MULTS_1_12(79)(PERCISION downto 1));
			MULTS_2_6(80)<=signed(MULTS_1_11(80)(PERCISION) & MULTS_1_11(80)(PERCISION downto 1))+signed(MULTS_1_12(80)(PERCISION) & MULTS_1_12(80)(PERCISION downto 1));
			MULTS_2_6(81)<=signed(MULTS_1_11(81)(PERCISION) & MULTS_1_11(81)(PERCISION downto 1))+signed(MULTS_1_12(81)(PERCISION) & MULTS_1_12(81)(PERCISION downto 1));
			MULTS_2_6(82)<=signed(MULTS_1_11(82)(PERCISION) & MULTS_1_11(82)(PERCISION downto 1))+signed(MULTS_1_12(82)(PERCISION) & MULTS_1_12(82)(PERCISION downto 1));
			MULTS_2_6(83)<=signed(MULTS_1_11(83)(PERCISION) & MULTS_1_11(83)(PERCISION downto 1))+signed(MULTS_1_12(83)(PERCISION) & MULTS_1_12(83)(PERCISION downto 1));

			MULTS_2_7(0)<=signed(MULTS_1_13(0)(PERCISION) & MULTS_1_13(0)(PERCISION downto 1))+signed(MULTS_1_14(0)(PERCISION) & MULTS_1_14(0)(PERCISION downto 1));
			MULTS_2_7(1)<=signed(MULTS_1_13(1)(PERCISION) & MULTS_1_13(1)(PERCISION downto 1))+signed(MULTS_1_14(1)(PERCISION) & MULTS_1_14(1)(PERCISION downto 1));
			MULTS_2_7(2)<=signed(MULTS_1_13(2)(PERCISION) & MULTS_1_13(2)(PERCISION downto 1))+signed(MULTS_1_14(2)(PERCISION) & MULTS_1_14(2)(PERCISION downto 1));
			MULTS_2_7(3)<=signed(MULTS_1_13(3)(PERCISION) & MULTS_1_13(3)(PERCISION downto 1))+signed(MULTS_1_14(3)(PERCISION) & MULTS_1_14(3)(PERCISION downto 1));
			MULTS_2_7(4)<=signed(MULTS_1_13(4)(PERCISION) & MULTS_1_13(4)(PERCISION downto 1))+signed(MULTS_1_14(4)(PERCISION) & MULTS_1_14(4)(PERCISION downto 1));
			MULTS_2_7(5)<=signed(MULTS_1_13(5)(PERCISION) & MULTS_1_13(5)(PERCISION downto 1))+signed(MULTS_1_14(5)(PERCISION) & MULTS_1_14(5)(PERCISION downto 1));
			MULTS_2_7(6)<=signed(MULTS_1_13(6)(PERCISION) & MULTS_1_13(6)(PERCISION downto 1))+signed(MULTS_1_14(6)(PERCISION) & MULTS_1_14(6)(PERCISION downto 1));
			MULTS_2_7(7)<=signed(MULTS_1_13(7)(PERCISION) & MULTS_1_13(7)(PERCISION downto 1))+signed(MULTS_1_14(7)(PERCISION) & MULTS_1_14(7)(PERCISION downto 1));
			MULTS_2_7(8)<=signed(MULTS_1_13(8)(PERCISION) & MULTS_1_13(8)(PERCISION downto 1))+signed(MULTS_1_14(8)(PERCISION) & MULTS_1_14(8)(PERCISION downto 1));
			MULTS_2_7(9)<=signed(MULTS_1_13(9)(PERCISION) & MULTS_1_13(9)(PERCISION downto 1))+signed(MULTS_1_14(9)(PERCISION) & MULTS_1_14(9)(PERCISION downto 1));
			MULTS_2_7(10)<=signed(MULTS_1_13(10)(PERCISION) & MULTS_1_13(10)(PERCISION downto 1))+signed(MULTS_1_14(10)(PERCISION) & MULTS_1_14(10)(PERCISION downto 1));
			MULTS_2_7(11)<=signed(MULTS_1_13(11)(PERCISION) & MULTS_1_13(11)(PERCISION downto 1))+signed(MULTS_1_14(11)(PERCISION) & MULTS_1_14(11)(PERCISION downto 1));
			MULTS_2_7(12)<=signed(MULTS_1_13(12)(PERCISION) & MULTS_1_13(12)(PERCISION downto 1))+signed(MULTS_1_14(12)(PERCISION) & MULTS_1_14(12)(PERCISION downto 1));
			MULTS_2_7(13)<=signed(MULTS_1_13(13)(PERCISION) & MULTS_1_13(13)(PERCISION downto 1))+signed(MULTS_1_14(13)(PERCISION) & MULTS_1_14(13)(PERCISION downto 1));
			MULTS_2_7(14)<=signed(MULTS_1_13(14)(PERCISION) & MULTS_1_13(14)(PERCISION downto 1))+signed(MULTS_1_14(14)(PERCISION) & MULTS_1_14(14)(PERCISION downto 1));
			MULTS_2_7(15)<=signed(MULTS_1_13(15)(PERCISION) & MULTS_1_13(15)(PERCISION downto 1))+signed(MULTS_1_14(15)(PERCISION) & MULTS_1_14(15)(PERCISION downto 1));
			MULTS_2_7(16)<=signed(MULTS_1_13(16)(PERCISION) & MULTS_1_13(16)(PERCISION downto 1))+signed(MULTS_1_14(16)(PERCISION) & MULTS_1_14(16)(PERCISION downto 1));
			MULTS_2_7(17)<=signed(MULTS_1_13(17)(PERCISION) & MULTS_1_13(17)(PERCISION downto 1))+signed(MULTS_1_14(17)(PERCISION) & MULTS_1_14(17)(PERCISION downto 1));
			MULTS_2_7(18)<=signed(MULTS_1_13(18)(PERCISION) & MULTS_1_13(18)(PERCISION downto 1))+signed(MULTS_1_14(18)(PERCISION) & MULTS_1_14(18)(PERCISION downto 1));
			MULTS_2_7(19)<=signed(MULTS_1_13(19)(PERCISION) & MULTS_1_13(19)(PERCISION downto 1))+signed(MULTS_1_14(19)(PERCISION) & MULTS_1_14(19)(PERCISION downto 1));
			MULTS_2_7(20)<=signed(MULTS_1_13(20)(PERCISION) & MULTS_1_13(20)(PERCISION downto 1))+signed(MULTS_1_14(20)(PERCISION) & MULTS_1_14(20)(PERCISION downto 1));
			MULTS_2_7(21)<=signed(MULTS_1_13(21)(PERCISION) & MULTS_1_13(21)(PERCISION downto 1))+signed(MULTS_1_14(21)(PERCISION) & MULTS_1_14(21)(PERCISION downto 1));
			MULTS_2_7(22)<=signed(MULTS_1_13(22)(PERCISION) & MULTS_1_13(22)(PERCISION downto 1))+signed(MULTS_1_14(22)(PERCISION) & MULTS_1_14(22)(PERCISION downto 1));
			MULTS_2_7(23)<=signed(MULTS_1_13(23)(PERCISION) & MULTS_1_13(23)(PERCISION downto 1))+signed(MULTS_1_14(23)(PERCISION) & MULTS_1_14(23)(PERCISION downto 1));
			MULTS_2_7(24)<=signed(MULTS_1_13(24)(PERCISION) & MULTS_1_13(24)(PERCISION downto 1))+signed(MULTS_1_14(24)(PERCISION) & MULTS_1_14(24)(PERCISION downto 1));
			MULTS_2_7(25)<=signed(MULTS_1_13(25)(PERCISION) & MULTS_1_13(25)(PERCISION downto 1))+signed(MULTS_1_14(25)(PERCISION) & MULTS_1_14(25)(PERCISION downto 1));
			MULTS_2_7(26)<=signed(MULTS_1_13(26)(PERCISION) & MULTS_1_13(26)(PERCISION downto 1))+signed(MULTS_1_14(26)(PERCISION) & MULTS_1_14(26)(PERCISION downto 1));
			MULTS_2_7(27)<=signed(MULTS_1_13(27)(PERCISION) & MULTS_1_13(27)(PERCISION downto 1))+signed(MULTS_1_14(27)(PERCISION) & MULTS_1_14(27)(PERCISION downto 1));
			MULTS_2_7(28)<=signed(MULTS_1_13(28)(PERCISION) & MULTS_1_13(28)(PERCISION downto 1))+signed(MULTS_1_14(28)(PERCISION) & MULTS_1_14(28)(PERCISION downto 1));
			MULTS_2_7(29)<=signed(MULTS_1_13(29)(PERCISION) & MULTS_1_13(29)(PERCISION downto 1))+signed(MULTS_1_14(29)(PERCISION) & MULTS_1_14(29)(PERCISION downto 1));
			MULTS_2_7(30)<=signed(MULTS_1_13(30)(PERCISION) & MULTS_1_13(30)(PERCISION downto 1))+signed(MULTS_1_14(30)(PERCISION) & MULTS_1_14(30)(PERCISION downto 1));
			MULTS_2_7(31)<=signed(MULTS_1_13(31)(PERCISION) & MULTS_1_13(31)(PERCISION downto 1))+signed(MULTS_1_14(31)(PERCISION) & MULTS_1_14(31)(PERCISION downto 1));
			MULTS_2_7(32)<=signed(MULTS_1_13(32)(PERCISION) & MULTS_1_13(32)(PERCISION downto 1))+signed(MULTS_1_14(32)(PERCISION) & MULTS_1_14(32)(PERCISION downto 1));
			MULTS_2_7(33)<=signed(MULTS_1_13(33)(PERCISION) & MULTS_1_13(33)(PERCISION downto 1))+signed(MULTS_1_14(33)(PERCISION) & MULTS_1_14(33)(PERCISION downto 1));
			MULTS_2_7(34)<=signed(MULTS_1_13(34)(PERCISION) & MULTS_1_13(34)(PERCISION downto 1))+signed(MULTS_1_14(34)(PERCISION) & MULTS_1_14(34)(PERCISION downto 1));
			MULTS_2_7(35)<=signed(MULTS_1_13(35)(PERCISION) & MULTS_1_13(35)(PERCISION downto 1))+signed(MULTS_1_14(35)(PERCISION) & MULTS_1_14(35)(PERCISION downto 1));
			MULTS_2_7(36)<=signed(MULTS_1_13(36)(PERCISION) & MULTS_1_13(36)(PERCISION downto 1))+signed(MULTS_1_14(36)(PERCISION) & MULTS_1_14(36)(PERCISION downto 1));
			MULTS_2_7(37)<=signed(MULTS_1_13(37)(PERCISION) & MULTS_1_13(37)(PERCISION downto 1))+signed(MULTS_1_14(37)(PERCISION) & MULTS_1_14(37)(PERCISION downto 1));
			MULTS_2_7(38)<=signed(MULTS_1_13(38)(PERCISION) & MULTS_1_13(38)(PERCISION downto 1))+signed(MULTS_1_14(38)(PERCISION) & MULTS_1_14(38)(PERCISION downto 1));
			MULTS_2_7(39)<=signed(MULTS_1_13(39)(PERCISION) & MULTS_1_13(39)(PERCISION downto 1))+signed(MULTS_1_14(39)(PERCISION) & MULTS_1_14(39)(PERCISION downto 1));
			MULTS_2_7(40)<=signed(MULTS_1_13(40)(PERCISION) & MULTS_1_13(40)(PERCISION downto 1))+signed(MULTS_1_14(40)(PERCISION) & MULTS_1_14(40)(PERCISION downto 1));
			MULTS_2_7(41)<=signed(MULTS_1_13(41)(PERCISION) & MULTS_1_13(41)(PERCISION downto 1))+signed(MULTS_1_14(41)(PERCISION) & MULTS_1_14(41)(PERCISION downto 1));
			MULTS_2_7(42)<=signed(MULTS_1_13(42)(PERCISION) & MULTS_1_13(42)(PERCISION downto 1))+signed(MULTS_1_14(42)(PERCISION) & MULTS_1_14(42)(PERCISION downto 1));
			MULTS_2_7(43)<=signed(MULTS_1_13(43)(PERCISION) & MULTS_1_13(43)(PERCISION downto 1))+signed(MULTS_1_14(43)(PERCISION) & MULTS_1_14(43)(PERCISION downto 1));
			MULTS_2_7(44)<=signed(MULTS_1_13(44)(PERCISION) & MULTS_1_13(44)(PERCISION downto 1))+signed(MULTS_1_14(44)(PERCISION) & MULTS_1_14(44)(PERCISION downto 1));
			MULTS_2_7(45)<=signed(MULTS_1_13(45)(PERCISION) & MULTS_1_13(45)(PERCISION downto 1))+signed(MULTS_1_14(45)(PERCISION) & MULTS_1_14(45)(PERCISION downto 1));
			MULTS_2_7(46)<=signed(MULTS_1_13(46)(PERCISION) & MULTS_1_13(46)(PERCISION downto 1))+signed(MULTS_1_14(46)(PERCISION) & MULTS_1_14(46)(PERCISION downto 1));
			MULTS_2_7(47)<=signed(MULTS_1_13(47)(PERCISION) & MULTS_1_13(47)(PERCISION downto 1))+signed(MULTS_1_14(47)(PERCISION) & MULTS_1_14(47)(PERCISION downto 1));
			MULTS_2_7(48)<=signed(MULTS_1_13(48)(PERCISION) & MULTS_1_13(48)(PERCISION downto 1))+signed(MULTS_1_14(48)(PERCISION) & MULTS_1_14(48)(PERCISION downto 1));
			MULTS_2_7(49)<=signed(MULTS_1_13(49)(PERCISION) & MULTS_1_13(49)(PERCISION downto 1))+signed(MULTS_1_14(49)(PERCISION) & MULTS_1_14(49)(PERCISION downto 1));
			MULTS_2_7(50)<=signed(MULTS_1_13(50)(PERCISION) & MULTS_1_13(50)(PERCISION downto 1))+signed(MULTS_1_14(50)(PERCISION) & MULTS_1_14(50)(PERCISION downto 1));
			MULTS_2_7(51)<=signed(MULTS_1_13(51)(PERCISION) & MULTS_1_13(51)(PERCISION downto 1))+signed(MULTS_1_14(51)(PERCISION) & MULTS_1_14(51)(PERCISION downto 1));
			MULTS_2_7(52)<=signed(MULTS_1_13(52)(PERCISION) & MULTS_1_13(52)(PERCISION downto 1))+signed(MULTS_1_14(52)(PERCISION) & MULTS_1_14(52)(PERCISION downto 1));
			MULTS_2_7(53)<=signed(MULTS_1_13(53)(PERCISION) & MULTS_1_13(53)(PERCISION downto 1))+signed(MULTS_1_14(53)(PERCISION) & MULTS_1_14(53)(PERCISION downto 1));
			MULTS_2_7(54)<=signed(MULTS_1_13(54)(PERCISION) & MULTS_1_13(54)(PERCISION downto 1))+signed(MULTS_1_14(54)(PERCISION) & MULTS_1_14(54)(PERCISION downto 1));
			MULTS_2_7(55)<=signed(MULTS_1_13(55)(PERCISION) & MULTS_1_13(55)(PERCISION downto 1))+signed(MULTS_1_14(55)(PERCISION) & MULTS_1_14(55)(PERCISION downto 1));
			MULTS_2_7(56)<=signed(MULTS_1_13(56)(PERCISION) & MULTS_1_13(56)(PERCISION downto 1))+signed(MULTS_1_14(56)(PERCISION) & MULTS_1_14(56)(PERCISION downto 1));
			MULTS_2_7(57)<=signed(MULTS_1_13(57)(PERCISION) & MULTS_1_13(57)(PERCISION downto 1))+signed(MULTS_1_14(57)(PERCISION) & MULTS_1_14(57)(PERCISION downto 1));
			MULTS_2_7(58)<=signed(MULTS_1_13(58)(PERCISION) & MULTS_1_13(58)(PERCISION downto 1))+signed(MULTS_1_14(58)(PERCISION) & MULTS_1_14(58)(PERCISION downto 1));
			MULTS_2_7(59)<=signed(MULTS_1_13(59)(PERCISION) & MULTS_1_13(59)(PERCISION downto 1))+signed(MULTS_1_14(59)(PERCISION) & MULTS_1_14(59)(PERCISION downto 1));
			MULTS_2_7(60)<=signed(MULTS_1_13(60)(PERCISION) & MULTS_1_13(60)(PERCISION downto 1))+signed(MULTS_1_14(60)(PERCISION) & MULTS_1_14(60)(PERCISION downto 1));
			MULTS_2_7(61)<=signed(MULTS_1_13(61)(PERCISION) & MULTS_1_13(61)(PERCISION downto 1))+signed(MULTS_1_14(61)(PERCISION) & MULTS_1_14(61)(PERCISION downto 1));
			MULTS_2_7(62)<=signed(MULTS_1_13(62)(PERCISION) & MULTS_1_13(62)(PERCISION downto 1))+signed(MULTS_1_14(62)(PERCISION) & MULTS_1_14(62)(PERCISION downto 1));
			MULTS_2_7(63)<=signed(MULTS_1_13(63)(PERCISION) & MULTS_1_13(63)(PERCISION downto 1))+signed(MULTS_1_14(63)(PERCISION) & MULTS_1_14(63)(PERCISION downto 1));
			MULTS_2_7(64)<=signed(MULTS_1_13(64)(PERCISION) & MULTS_1_13(64)(PERCISION downto 1))+signed(MULTS_1_14(64)(PERCISION) & MULTS_1_14(64)(PERCISION downto 1));
			MULTS_2_7(65)<=signed(MULTS_1_13(65)(PERCISION) & MULTS_1_13(65)(PERCISION downto 1))+signed(MULTS_1_14(65)(PERCISION) & MULTS_1_14(65)(PERCISION downto 1));
			MULTS_2_7(66)<=signed(MULTS_1_13(66)(PERCISION) & MULTS_1_13(66)(PERCISION downto 1))+signed(MULTS_1_14(66)(PERCISION) & MULTS_1_14(66)(PERCISION downto 1));
			MULTS_2_7(67)<=signed(MULTS_1_13(67)(PERCISION) & MULTS_1_13(67)(PERCISION downto 1))+signed(MULTS_1_14(67)(PERCISION) & MULTS_1_14(67)(PERCISION downto 1));
			MULTS_2_7(68)<=signed(MULTS_1_13(68)(PERCISION) & MULTS_1_13(68)(PERCISION downto 1))+signed(MULTS_1_14(68)(PERCISION) & MULTS_1_14(68)(PERCISION downto 1));
			MULTS_2_7(69)<=signed(MULTS_1_13(69)(PERCISION) & MULTS_1_13(69)(PERCISION downto 1))+signed(MULTS_1_14(69)(PERCISION) & MULTS_1_14(69)(PERCISION downto 1));
			MULTS_2_7(70)<=signed(MULTS_1_13(70)(PERCISION) & MULTS_1_13(70)(PERCISION downto 1))+signed(MULTS_1_14(70)(PERCISION) & MULTS_1_14(70)(PERCISION downto 1));
			MULTS_2_7(71)<=signed(MULTS_1_13(71)(PERCISION) & MULTS_1_13(71)(PERCISION downto 1))+signed(MULTS_1_14(71)(PERCISION) & MULTS_1_14(71)(PERCISION downto 1));
			MULTS_2_7(72)<=signed(MULTS_1_13(72)(PERCISION) & MULTS_1_13(72)(PERCISION downto 1))+signed(MULTS_1_14(72)(PERCISION) & MULTS_1_14(72)(PERCISION downto 1));
			MULTS_2_7(73)<=signed(MULTS_1_13(73)(PERCISION) & MULTS_1_13(73)(PERCISION downto 1))+signed(MULTS_1_14(73)(PERCISION) & MULTS_1_14(73)(PERCISION downto 1));
			MULTS_2_7(74)<=signed(MULTS_1_13(74)(PERCISION) & MULTS_1_13(74)(PERCISION downto 1))+signed(MULTS_1_14(74)(PERCISION) & MULTS_1_14(74)(PERCISION downto 1));
			MULTS_2_7(75)<=signed(MULTS_1_13(75)(PERCISION) & MULTS_1_13(75)(PERCISION downto 1))+signed(MULTS_1_14(75)(PERCISION) & MULTS_1_14(75)(PERCISION downto 1));
			MULTS_2_7(76)<=signed(MULTS_1_13(76)(PERCISION) & MULTS_1_13(76)(PERCISION downto 1))+signed(MULTS_1_14(76)(PERCISION) & MULTS_1_14(76)(PERCISION downto 1));
			MULTS_2_7(77)<=signed(MULTS_1_13(77)(PERCISION) & MULTS_1_13(77)(PERCISION downto 1))+signed(MULTS_1_14(77)(PERCISION) & MULTS_1_14(77)(PERCISION downto 1));
			MULTS_2_7(78)<=signed(MULTS_1_13(78)(PERCISION) & MULTS_1_13(78)(PERCISION downto 1))+signed(MULTS_1_14(78)(PERCISION) & MULTS_1_14(78)(PERCISION downto 1));
			MULTS_2_7(79)<=signed(MULTS_1_13(79)(PERCISION) & MULTS_1_13(79)(PERCISION downto 1))+signed(MULTS_1_14(79)(PERCISION) & MULTS_1_14(79)(PERCISION downto 1));
			MULTS_2_7(80)<=signed(MULTS_1_13(80)(PERCISION) & MULTS_1_13(80)(PERCISION downto 1))+signed(MULTS_1_14(80)(PERCISION) & MULTS_1_14(80)(PERCISION downto 1));
			MULTS_2_7(81)<=signed(MULTS_1_13(81)(PERCISION) & MULTS_1_13(81)(PERCISION downto 1))+signed(MULTS_1_14(81)(PERCISION) & MULTS_1_14(81)(PERCISION downto 1));
			MULTS_2_7(82)<=signed(MULTS_1_13(82)(PERCISION) & MULTS_1_13(82)(PERCISION downto 1))+signed(MULTS_1_14(82)(PERCISION) & MULTS_1_14(82)(PERCISION downto 1));
			MULTS_2_7(83)<=signed(MULTS_1_13(83)(PERCISION) & MULTS_1_13(83)(PERCISION downto 1))+signed(MULTS_1_14(83)(PERCISION) & MULTS_1_14(83)(PERCISION downto 1));

			MULTS_2_8(0)<=signed(MULTS_1_15(0)(PERCISION) & MULTS_1_15(0)(PERCISION downto 1))+signed(MULTS_1_16(0)(PERCISION) & MULTS_1_16(0)(PERCISION downto 1));
			MULTS_2_8(1)<=signed(MULTS_1_15(1)(PERCISION) & MULTS_1_15(1)(PERCISION downto 1))+signed(MULTS_1_16(1)(PERCISION) & MULTS_1_16(1)(PERCISION downto 1));
			MULTS_2_8(2)<=signed(MULTS_1_15(2)(PERCISION) & MULTS_1_15(2)(PERCISION downto 1))+signed(MULTS_1_16(2)(PERCISION) & MULTS_1_16(2)(PERCISION downto 1));
			MULTS_2_8(3)<=signed(MULTS_1_15(3)(PERCISION) & MULTS_1_15(3)(PERCISION downto 1))+signed(MULTS_1_16(3)(PERCISION) & MULTS_1_16(3)(PERCISION downto 1));
			MULTS_2_8(4)<=signed(MULTS_1_15(4)(PERCISION) & MULTS_1_15(4)(PERCISION downto 1))+signed(MULTS_1_16(4)(PERCISION) & MULTS_1_16(4)(PERCISION downto 1));
			MULTS_2_8(5)<=signed(MULTS_1_15(5)(PERCISION) & MULTS_1_15(5)(PERCISION downto 1))+signed(MULTS_1_16(5)(PERCISION) & MULTS_1_16(5)(PERCISION downto 1));
			MULTS_2_8(6)<=signed(MULTS_1_15(6)(PERCISION) & MULTS_1_15(6)(PERCISION downto 1))+signed(MULTS_1_16(6)(PERCISION) & MULTS_1_16(6)(PERCISION downto 1));
			MULTS_2_8(7)<=signed(MULTS_1_15(7)(PERCISION) & MULTS_1_15(7)(PERCISION downto 1))+signed(MULTS_1_16(7)(PERCISION) & MULTS_1_16(7)(PERCISION downto 1));
			MULTS_2_8(8)<=signed(MULTS_1_15(8)(PERCISION) & MULTS_1_15(8)(PERCISION downto 1))+signed(MULTS_1_16(8)(PERCISION) & MULTS_1_16(8)(PERCISION downto 1));
			MULTS_2_8(9)<=signed(MULTS_1_15(9)(PERCISION) & MULTS_1_15(9)(PERCISION downto 1))+signed(MULTS_1_16(9)(PERCISION) & MULTS_1_16(9)(PERCISION downto 1));
			MULTS_2_8(10)<=signed(MULTS_1_15(10)(PERCISION) & MULTS_1_15(10)(PERCISION downto 1))+signed(MULTS_1_16(10)(PERCISION) & MULTS_1_16(10)(PERCISION downto 1));
			MULTS_2_8(11)<=signed(MULTS_1_15(11)(PERCISION) & MULTS_1_15(11)(PERCISION downto 1))+signed(MULTS_1_16(11)(PERCISION) & MULTS_1_16(11)(PERCISION downto 1));
			MULTS_2_8(12)<=signed(MULTS_1_15(12)(PERCISION) & MULTS_1_15(12)(PERCISION downto 1))+signed(MULTS_1_16(12)(PERCISION) & MULTS_1_16(12)(PERCISION downto 1));
			MULTS_2_8(13)<=signed(MULTS_1_15(13)(PERCISION) & MULTS_1_15(13)(PERCISION downto 1))+signed(MULTS_1_16(13)(PERCISION) & MULTS_1_16(13)(PERCISION downto 1));
			MULTS_2_8(14)<=signed(MULTS_1_15(14)(PERCISION) & MULTS_1_15(14)(PERCISION downto 1))+signed(MULTS_1_16(14)(PERCISION) & MULTS_1_16(14)(PERCISION downto 1));
			MULTS_2_8(15)<=signed(MULTS_1_15(15)(PERCISION) & MULTS_1_15(15)(PERCISION downto 1))+signed(MULTS_1_16(15)(PERCISION) & MULTS_1_16(15)(PERCISION downto 1));
			MULTS_2_8(16)<=signed(MULTS_1_15(16)(PERCISION) & MULTS_1_15(16)(PERCISION downto 1))+signed(MULTS_1_16(16)(PERCISION) & MULTS_1_16(16)(PERCISION downto 1));
			MULTS_2_8(17)<=signed(MULTS_1_15(17)(PERCISION) & MULTS_1_15(17)(PERCISION downto 1))+signed(MULTS_1_16(17)(PERCISION) & MULTS_1_16(17)(PERCISION downto 1));
			MULTS_2_8(18)<=signed(MULTS_1_15(18)(PERCISION) & MULTS_1_15(18)(PERCISION downto 1))+signed(MULTS_1_16(18)(PERCISION) & MULTS_1_16(18)(PERCISION downto 1));
			MULTS_2_8(19)<=signed(MULTS_1_15(19)(PERCISION) & MULTS_1_15(19)(PERCISION downto 1))+signed(MULTS_1_16(19)(PERCISION) & MULTS_1_16(19)(PERCISION downto 1));
			MULTS_2_8(20)<=signed(MULTS_1_15(20)(PERCISION) & MULTS_1_15(20)(PERCISION downto 1))+signed(MULTS_1_16(20)(PERCISION) & MULTS_1_16(20)(PERCISION downto 1));
			MULTS_2_8(21)<=signed(MULTS_1_15(21)(PERCISION) & MULTS_1_15(21)(PERCISION downto 1))+signed(MULTS_1_16(21)(PERCISION) & MULTS_1_16(21)(PERCISION downto 1));
			MULTS_2_8(22)<=signed(MULTS_1_15(22)(PERCISION) & MULTS_1_15(22)(PERCISION downto 1))+signed(MULTS_1_16(22)(PERCISION) & MULTS_1_16(22)(PERCISION downto 1));
			MULTS_2_8(23)<=signed(MULTS_1_15(23)(PERCISION) & MULTS_1_15(23)(PERCISION downto 1))+signed(MULTS_1_16(23)(PERCISION) & MULTS_1_16(23)(PERCISION downto 1));
			MULTS_2_8(24)<=signed(MULTS_1_15(24)(PERCISION) & MULTS_1_15(24)(PERCISION downto 1))+signed(MULTS_1_16(24)(PERCISION) & MULTS_1_16(24)(PERCISION downto 1));
			MULTS_2_8(25)<=signed(MULTS_1_15(25)(PERCISION) & MULTS_1_15(25)(PERCISION downto 1))+signed(MULTS_1_16(25)(PERCISION) & MULTS_1_16(25)(PERCISION downto 1));
			MULTS_2_8(26)<=signed(MULTS_1_15(26)(PERCISION) & MULTS_1_15(26)(PERCISION downto 1))+signed(MULTS_1_16(26)(PERCISION) & MULTS_1_16(26)(PERCISION downto 1));
			MULTS_2_8(27)<=signed(MULTS_1_15(27)(PERCISION) & MULTS_1_15(27)(PERCISION downto 1))+signed(MULTS_1_16(27)(PERCISION) & MULTS_1_16(27)(PERCISION downto 1));
			MULTS_2_8(28)<=signed(MULTS_1_15(28)(PERCISION) & MULTS_1_15(28)(PERCISION downto 1))+signed(MULTS_1_16(28)(PERCISION) & MULTS_1_16(28)(PERCISION downto 1));
			MULTS_2_8(29)<=signed(MULTS_1_15(29)(PERCISION) & MULTS_1_15(29)(PERCISION downto 1))+signed(MULTS_1_16(29)(PERCISION) & MULTS_1_16(29)(PERCISION downto 1));
			MULTS_2_8(30)<=signed(MULTS_1_15(30)(PERCISION) & MULTS_1_15(30)(PERCISION downto 1))+signed(MULTS_1_16(30)(PERCISION) & MULTS_1_16(30)(PERCISION downto 1));
			MULTS_2_8(31)<=signed(MULTS_1_15(31)(PERCISION) & MULTS_1_15(31)(PERCISION downto 1))+signed(MULTS_1_16(31)(PERCISION) & MULTS_1_16(31)(PERCISION downto 1));
			MULTS_2_8(32)<=signed(MULTS_1_15(32)(PERCISION) & MULTS_1_15(32)(PERCISION downto 1))+signed(MULTS_1_16(32)(PERCISION) & MULTS_1_16(32)(PERCISION downto 1));
			MULTS_2_8(33)<=signed(MULTS_1_15(33)(PERCISION) & MULTS_1_15(33)(PERCISION downto 1))+signed(MULTS_1_16(33)(PERCISION) & MULTS_1_16(33)(PERCISION downto 1));
			MULTS_2_8(34)<=signed(MULTS_1_15(34)(PERCISION) & MULTS_1_15(34)(PERCISION downto 1))+signed(MULTS_1_16(34)(PERCISION) & MULTS_1_16(34)(PERCISION downto 1));
			MULTS_2_8(35)<=signed(MULTS_1_15(35)(PERCISION) & MULTS_1_15(35)(PERCISION downto 1))+signed(MULTS_1_16(35)(PERCISION) & MULTS_1_16(35)(PERCISION downto 1));
			MULTS_2_8(36)<=signed(MULTS_1_15(36)(PERCISION) & MULTS_1_15(36)(PERCISION downto 1))+signed(MULTS_1_16(36)(PERCISION) & MULTS_1_16(36)(PERCISION downto 1));
			MULTS_2_8(37)<=signed(MULTS_1_15(37)(PERCISION) & MULTS_1_15(37)(PERCISION downto 1))+signed(MULTS_1_16(37)(PERCISION) & MULTS_1_16(37)(PERCISION downto 1));
			MULTS_2_8(38)<=signed(MULTS_1_15(38)(PERCISION) & MULTS_1_15(38)(PERCISION downto 1))+signed(MULTS_1_16(38)(PERCISION) & MULTS_1_16(38)(PERCISION downto 1));
			MULTS_2_8(39)<=signed(MULTS_1_15(39)(PERCISION) & MULTS_1_15(39)(PERCISION downto 1))+signed(MULTS_1_16(39)(PERCISION) & MULTS_1_16(39)(PERCISION downto 1));
			MULTS_2_8(40)<=signed(MULTS_1_15(40)(PERCISION) & MULTS_1_15(40)(PERCISION downto 1))+signed(MULTS_1_16(40)(PERCISION) & MULTS_1_16(40)(PERCISION downto 1));
			MULTS_2_8(41)<=signed(MULTS_1_15(41)(PERCISION) & MULTS_1_15(41)(PERCISION downto 1))+signed(MULTS_1_16(41)(PERCISION) & MULTS_1_16(41)(PERCISION downto 1));
			MULTS_2_8(42)<=signed(MULTS_1_15(42)(PERCISION) & MULTS_1_15(42)(PERCISION downto 1))+signed(MULTS_1_16(42)(PERCISION) & MULTS_1_16(42)(PERCISION downto 1));
			MULTS_2_8(43)<=signed(MULTS_1_15(43)(PERCISION) & MULTS_1_15(43)(PERCISION downto 1))+signed(MULTS_1_16(43)(PERCISION) & MULTS_1_16(43)(PERCISION downto 1));
			MULTS_2_8(44)<=signed(MULTS_1_15(44)(PERCISION) & MULTS_1_15(44)(PERCISION downto 1))+signed(MULTS_1_16(44)(PERCISION) & MULTS_1_16(44)(PERCISION downto 1));
			MULTS_2_8(45)<=signed(MULTS_1_15(45)(PERCISION) & MULTS_1_15(45)(PERCISION downto 1))+signed(MULTS_1_16(45)(PERCISION) & MULTS_1_16(45)(PERCISION downto 1));
			MULTS_2_8(46)<=signed(MULTS_1_15(46)(PERCISION) & MULTS_1_15(46)(PERCISION downto 1))+signed(MULTS_1_16(46)(PERCISION) & MULTS_1_16(46)(PERCISION downto 1));
			MULTS_2_8(47)<=signed(MULTS_1_15(47)(PERCISION) & MULTS_1_15(47)(PERCISION downto 1))+signed(MULTS_1_16(47)(PERCISION) & MULTS_1_16(47)(PERCISION downto 1));
			MULTS_2_8(48)<=signed(MULTS_1_15(48)(PERCISION) & MULTS_1_15(48)(PERCISION downto 1))+signed(MULTS_1_16(48)(PERCISION) & MULTS_1_16(48)(PERCISION downto 1));
			MULTS_2_8(49)<=signed(MULTS_1_15(49)(PERCISION) & MULTS_1_15(49)(PERCISION downto 1))+signed(MULTS_1_16(49)(PERCISION) & MULTS_1_16(49)(PERCISION downto 1));
			MULTS_2_8(50)<=signed(MULTS_1_15(50)(PERCISION) & MULTS_1_15(50)(PERCISION downto 1))+signed(MULTS_1_16(50)(PERCISION) & MULTS_1_16(50)(PERCISION downto 1));
			MULTS_2_8(51)<=signed(MULTS_1_15(51)(PERCISION) & MULTS_1_15(51)(PERCISION downto 1))+signed(MULTS_1_16(51)(PERCISION) & MULTS_1_16(51)(PERCISION downto 1));
			MULTS_2_8(52)<=signed(MULTS_1_15(52)(PERCISION) & MULTS_1_15(52)(PERCISION downto 1))+signed(MULTS_1_16(52)(PERCISION) & MULTS_1_16(52)(PERCISION downto 1));
			MULTS_2_8(53)<=signed(MULTS_1_15(53)(PERCISION) & MULTS_1_15(53)(PERCISION downto 1))+signed(MULTS_1_16(53)(PERCISION) & MULTS_1_16(53)(PERCISION downto 1));
			MULTS_2_8(54)<=signed(MULTS_1_15(54)(PERCISION) & MULTS_1_15(54)(PERCISION downto 1))+signed(MULTS_1_16(54)(PERCISION) & MULTS_1_16(54)(PERCISION downto 1));
			MULTS_2_8(55)<=signed(MULTS_1_15(55)(PERCISION) & MULTS_1_15(55)(PERCISION downto 1))+signed(MULTS_1_16(55)(PERCISION) & MULTS_1_16(55)(PERCISION downto 1));
			MULTS_2_8(56)<=signed(MULTS_1_15(56)(PERCISION) & MULTS_1_15(56)(PERCISION downto 1))+signed(MULTS_1_16(56)(PERCISION) & MULTS_1_16(56)(PERCISION downto 1));
			MULTS_2_8(57)<=signed(MULTS_1_15(57)(PERCISION) & MULTS_1_15(57)(PERCISION downto 1))+signed(MULTS_1_16(57)(PERCISION) & MULTS_1_16(57)(PERCISION downto 1));
			MULTS_2_8(58)<=signed(MULTS_1_15(58)(PERCISION) & MULTS_1_15(58)(PERCISION downto 1))+signed(MULTS_1_16(58)(PERCISION) & MULTS_1_16(58)(PERCISION downto 1));
			MULTS_2_8(59)<=signed(MULTS_1_15(59)(PERCISION) & MULTS_1_15(59)(PERCISION downto 1))+signed(MULTS_1_16(59)(PERCISION) & MULTS_1_16(59)(PERCISION downto 1));
			MULTS_2_8(60)<=signed(MULTS_1_15(60)(PERCISION) & MULTS_1_15(60)(PERCISION downto 1))+signed(MULTS_1_16(60)(PERCISION) & MULTS_1_16(60)(PERCISION downto 1));
			MULTS_2_8(61)<=signed(MULTS_1_15(61)(PERCISION) & MULTS_1_15(61)(PERCISION downto 1))+signed(MULTS_1_16(61)(PERCISION) & MULTS_1_16(61)(PERCISION downto 1));
			MULTS_2_8(62)<=signed(MULTS_1_15(62)(PERCISION) & MULTS_1_15(62)(PERCISION downto 1))+signed(MULTS_1_16(62)(PERCISION) & MULTS_1_16(62)(PERCISION downto 1));
			MULTS_2_8(63)<=signed(MULTS_1_15(63)(PERCISION) & MULTS_1_15(63)(PERCISION downto 1))+signed(MULTS_1_16(63)(PERCISION) & MULTS_1_16(63)(PERCISION downto 1));
			MULTS_2_8(64)<=signed(MULTS_1_15(64)(PERCISION) & MULTS_1_15(64)(PERCISION downto 1))+signed(MULTS_1_16(64)(PERCISION) & MULTS_1_16(64)(PERCISION downto 1));
			MULTS_2_8(65)<=signed(MULTS_1_15(65)(PERCISION) & MULTS_1_15(65)(PERCISION downto 1))+signed(MULTS_1_16(65)(PERCISION) & MULTS_1_16(65)(PERCISION downto 1));
			MULTS_2_8(66)<=signed(MULTS_1_15(66)(PERCISION) & MULTS_1_15(66)(PERCISION downto 1))+signed(MULTS_1_16(66)(PERCISION) & MULTS_1_16(66)(PERCISION downto 1));
			MULTS_2_8(67)<=signed(MULTS_1_15(67)(PERCISION) & MULTS_1_15(67)(PERCISION downto 1))+signed(MULTS_1_16(67)(PERCISION) & MULTS_1_16(67)(PERCISION downto 1));
			MULTS_2_8(68)<=signed(MULTS_1_15(68)(PERCISION) & MULTS_1_15(68)(PERCISION downto 1))+signed(MULTS_1_16(68)(PERCISION) & MULTS_1_16(68)(PERCISION downto 1));
			MULTS_2_8(69)<=signed(MULTS_1_15(69)(PERCISION) & MULTS_1_15(69)(PERCISION downto 1))+signed(MULTS_1_16(69)(PERCISION) & MULTS_1_16(69)(PERCISION downto 1));
			MULTS_2_8(70)<=signed(MULTS_1_15(70)(PERCISION) & MULTS_1_15(70)(PERCISION downto 1))+signed(MULTS_1_16(70)(PERCISION) & MULTS_1_16(70)(PERCISION downto 1));
			MULTS_2_8(71)<=signed(MULTS_1_15(71)(PERCISION) & MULTS_1_15(71)(PERCISION downto 1))+signed(MULTS_1_16(71)(PERCISION) & MULTS_1_16(71)(PERCISION downto 1));
			MULTS_2_8(72)<=signed(MULTS_1_15(72)(PERCISION) & MULTS_1_15(72)(PERCISION downto 1))+signed(MULTS_1_16(72)(PERCISION) & MULTS_1_16(72)(PERCISION downto 1));
			MULTS_2_8(73)<=signed(MULTS_1_15(73)(PERCISION) & MULTS_1_15(73)(PERCISION downto 1))+signed(MULTS_1_16(73)(PERCISION) & MULTS_1_16(73)(PERCISION downto 1));
			MULTS_2_8(74)<=signed(MULTS_1_15(74)(PERCISION) & MULTS_1_15(74)(PERCISION downto 1))+signed(MULTS_1_16(74)(PERCISION) & MULTS_1_16(74)(PERCISION downto 1));
			MULTS_2_8(75)<=signed(MULTS_1_15(75)(PERCISION) & MULTS_1_15(75)(PERCISION downto 1))+signed(MULTS_1_16(75)(PERCISION) & MULTS_1_16(75)(PERCISION downto 1));
			MULTS_2_8(76)<=signed(MULTS_1_15(76)(PERCISION) & MULTS_1_15(76)(PERCISION downto 1))+signed(MULTS_1_16(76)(PERCISION) & MULTS_1_16(76)(PERCISION downto 1));
			MULTS_2_8(77)<=signed(MULTS_1_15(77)(PERCISION) & MULTS_1_15(77)(PERCISION downto 1))+signed(MULTS_1_16(77)(PERCISION) & MULTS_1_16(77)(PERCISION downto 1));
			MULTS_2_8(78)<=signed(MULTS_1_15(78)(PERCISION) & MULTS_1_15(78)(PERCISION downto 1))+signed(MULTS_1_16(78)(PERCISION) & MULTS_1_16(78)(PERCISION downto 1));
			MULTS_2_8(79)<=signed(MULTS_1_15(79)(PERCISION) & MULTS_1_15(79)(PERCISION downto 1))+signed(MULTS_1_16(79)(PERCISION) & MULTS_1_16(79)(PERCISION downto 1));
			MULTS_2_8(80)<=signed(MULTS_1_15(80)(PERCISION) & MULTS_1_15(80)(PERCISION downto 1))+signed(MULTS_1_16(80)(PERCISION) & MULTS_1_16(80)(PERCISION downto 1));
			MULTS_2_8(81)<=signed(MULTS_1_15(81)(PERCISION) & MULTS_1_15(81)(PERCISION downto 1))+signed(MULTS_1_16(81)(PERCISION) & MULTS_1_16(81)(PERCISION downto 1));
			MULTS_2_8(82)<=signed(MULTS_1_15(82)(PERCISION) & MULTS_1_15(82)(PERCISION downto 1))+signed(MULTS_1_16(82)(PERCISION) & MULTS_1_16(82)(PERCISION downto 1));
			MULTS_2_8(83)<=signed(MULTS_1_15(83)(PERCISION) & MULTS_1_15(83)(PERCISION downto 1))+signed(MULTS_1_16(83)(PERCISION) & MULTS_1_16(83)(PERCISION downto 1));

			MULTS_2_9(0)<=signed(MULTS_1_17(0)(PERCISION) & MULTS_1_17(0)(PERCISION downto 1))+signed(MULTS_1_18(0)(PERCISION) & MULTS_1_18(0)(PERCISION downto 1));
			MULTS_2_9(1)<=signed(MULTS_1_17(1)(PERCISION) & MULTS_1_17(1)(PERCISION downto 1))+signed(MULTS_1_18(1)(PERCISION) & MULTS_1_18(1)(PERCISION downto 1));
			MULTS_2_9(2)<=signed(MULTS_1_17(2)(PERCISION) & MULTS_1_17(2)(PERCISION downto 1))+signed(MULTS_1_18(2)(PERCISION) & MULTS_1_18(2)(PERCISION downto 1));
			MULTS_2_9(3)<=signed(MULTS_1_17(3)(PERCISION) & MULTS_1_17(3)(PERCISION downto 1))+signed(MULTS_1_18(3)(PERCISION) & MULTS_1_18(3)(PERCISION downto 1));
			MULTS_2_9(4)<=signed(MULTS_1_17(4)(PERCISION) & MULTS_1_17(4)(PERCISION downto 1))+signed(MULTS_1_18(4)(PERCISION) & MULTS_1_18(4)(PERCISION downto 1));
			MULTS_2_9(5)<=signed(MULTS_1_17(5)(PERCISION) & MULTS_1_17(5)(PERCISION downto 1))+signed(MULTS_1_18(5)(PERCISION) & MULTS_1_18(5)(PERCISION downto 1));
			MULTS_2_9(6)<=signed(MULTS_1_17(6)(PERCISION) & MULTS_1_17(6)(PERCISION downto 1))+signed(MULTS_1_18(6)(PERCISION) & MULTS_1_18(6)(PERCISION downto 1));
			MULTS_2_9(7)<=signed(MULTS_1_17(7)(PERCISION) & MULTS_1_17(7)(PERCISION downto 1))+signed(MULTS_1_18(7)(PERCISION) & MULTS_1_18(7)(PERCISION downto 1));
			MULTS_2_9(8)<=signed(MULTS_1_17(8)(PERCISION) & MULTS_1_17(8)(PERCISION downto 1))+signed(MULTS_1_18(8)(PERCISION) & MULTS_1_18(8)(PERCISION downto 1));
			MULTS_2_9(9)<=signed(MULTS_1_17(9)(PERCISION) & MULTS_1_17(9)(PERCISION downto 1))+signed(MULTS_1_18(9)(PERCISION) & MULTS_1_18(9)(PERCISION downto 1));
			MULTS_2_9(10)<=signed(MULTS_1_17(10)(PERCISION) & MULTS_1_17(10)(PERCISION downto 1))+signed(MULTS_1_18(10)(PERCISION) & MULTS_1_18(10)(PERCISION downto 1));
			MULTS_2_9(11)<=signed(MULTS_1_17(11)(PERCISION) & MULTS_1_17(11)(PERCISION downto 1))+signed(MULTS_1_18(11)(PERCISION) & MULTS_1_18(11)(PERCISION downto 1));
			MULTS_2_9(12)<=signed(MULTS_1_17(12)(PERCISION) & MULTS_1_17(12)(PERCISION downto 1))+signed(MULTS_1_18(12)(PERCISION) & MULTS_1_18(12)(PERCISION downto 1));
			MULTS_2_9(13)<=signed(MULTS_1_17(13)(PERCISION) & MULTS_1_17(13)(PERCISION downto 1))+signed(MULTS_1_18(13)(PERCISION) & MULTS_1_18(13)(PERCISION downto 1));
			MULTS_2_9(14)<=signed(MULTS_1_17(14)(PERCISION) & MULTS_1_17(14)(PERCISION downto 1))+signed(MULTS_1_18(14)(PERCISION) & MULTS_1_18(14)(PERCISION downto 1));
			MULTS_2_9(15)<=signed(MULTS_1_17(15)(PERCISION) & MULTS_1_17(15)(PERCISION downto 1))+signed(MULTS_1_18(15)(PERCISION) & MULTS_1_18(15)(PERCISION downto 1));
			MULTS_2_9(16)<=signed(MULTS_1_17(16)(PERCISION) & MULTS_1_17(16)(PERCISION downto 1))+signed(MULTS_1_18(16)(PERCISION) & MULTS_1_18(16)(PERCISION downto 1));
			MULTS_2_9(17)<=signed(MULTS_1_17(17)(PERCISION) & MULTS_1_17(17)(PERCISION downto 1))+signed(MULTS_1_18(17)(PERCISION) & MULTS_1_18(17)(PERCISION downto 1));
			MULTS_2_9(18)<=signed(MULTS_1_17(18)(PERCISION) & MULTS_1_17(18)(PERCISION downto 1))+signed(MULTS_1_18(18)(PERCISION) & MULTS_1_18(18)(PERCISION downto 1));
			MULTS_2_9(19)<=signed(MULTS_1_17(19)(PERCISION) & MULTS_1_17(19)(PERCISION downto 1))+signed(MULTS_1_18(19)(PERCISION) & MULTS_1_18(19)(PERCISION downto 1));
			MULTS_2_9(20)<=signed(MULTS_1_17(20)(PERCISION) & MULTS_1_17(20)(PERCISION downto 1))+signed(MULTS_1_18(20)(PERCISION) & MULTS_1_18(20)(PERCISION downto 1));
			MULTS_2_9(21)<=signed(MULTS_1_17(21)(PERCISION) & MULTS_1_17(21)(PERCISION downto 1))+signed(MULTS_1_18(21)(PERCISION) & MULTS_1_18(21)(PERCISION downto 1));
			MULTS_2_9(22)<=signed(MULTS_1_17(22)(PERCISION) & MULTS_1_17(22)(PERCISION downto 1))+signed(MULTS_1_18(22)(PERCISION) & MULTS_1_18(22)(PERCISION downto 1));
			MULTS_2_9(23)<=signed(MULTS_1_17(23)(PERCISION) & MULTS_1_17(23)(PERCISION downto 1))+signed(MULTS_1_18(23)(PERCISION) & MULTS_1_18(23)(PERCISION downto 1));
			MULTS_2_9(24)<=signed(MULTS_1_17(24)(PERCISION) & MULTS_1_17(24)(PERCISION downto 1))+signed(MULTS_1_18(24)(PERCISION) & MULTS_1_18(24)(PERCISION downto 1));
			MULTS_2_9(25)<=signed(MULTS_1_17(25)(PERCISION) & MULTS_1_17(25)(PERCISION downto 1))+signed(MULTS_1_18(25)(PERCISION) & MULTS_1_18(25)(PERCISION downto 1));
			MULTS_2_9(26)<=signed(MULTS_1_17(26)(PERCISION) & MULTS_1_17(26)(PERCISION downto 1))+signed(MULTS_1_18(26)(PERCISION) & MULTS_1_18(26)(PERCISION downto 1));
			MULTS_2_9(27)<=signed(MULTS_1_17(27)(PERCISION) & MULTS_1_17(27)(PERCISION downto 1))+signed(MULTS_1_18(27)(PERCISION) & MULTS_1_18(27)(PERCISION downto 1));
			MULTS_2_9(28)<=signed(MULTS_1_17(28)(PERCISION) & MULTS_1_17(28)(PERCISION downto 1))+signed(MULTS_1_18(28)(PERCISION) & MULTS_1_18(28)(PERCISION downto 1));
			MULTS_2_9(29)<=signed(MULTS_1_17(29)(PERCISION) & MULTS_1_17(29)(PERCISION downto 1))+signed(MULTS_1_18(29)(PERCISION) & MULTS_1_18(29)(PERCISION downto 1));
			MULTS_2_9(30)<=signed(MULTS_1_17(30)(PERCISION) & MULTS_1_17(30)(PERCISION downto 1))+signed(MULTS_1_18(30)(PERCISION) & MULTS_1_18(30)(PERCISION downto 1));
			MULTS_2_9(31)<=signed(MULTS_1_17(31)(PERCISION) & MULTS_1_17(31)(PERCISION downto 1))+signed(MULTS_1_18(31)(PERCISION) & MULTS_1_18(31)(PERCISION downto 1));
			MULTS_2_9(32)<=signed(MULTS_1_17(32)(PERCISION) & MULTS_1_17(32)(PERCISION downto 1))+signed(MULTS_1_18(32)(PERCISION) & MULTS_1_18(32)(PERCISION downto 1));
			MULTS_2_9(33)<=signed(MULTS_1_17(33)(PERCISION) & MULTS_1_17(33)(PERCISION downto 1))+signed(MULTS_1_18(33)(PERCISION) & MULTS_1_18(33)(PERCISION downto 1));
			MULTS_2_9(34)<=signed(MULTS_1_17(34)(PERCISION) & MULTS_1_17(34)(PERCISION downto 1))+signed(MULTS_1_18(34)(PERCISION) & MULTS_1_18(34)(PERCISION downto 1));
			MULTS_2_9(35)<=signed(MULTS_1_17(35)(PERCISION) & MULTS_1_17(35)(PERCISION downto 1))+signed(MULTS_1_18(35)(PERCISION) & MULTS_1_18(35)(PERCISION downto 1));
			MULTS_2_9(36)<=signed(MULTS_1_17(36)(PERCISION) & MULTS_1_17(36)(PERCISION downto 1))+signed(MULTS_1_18(36)(PERCISION) & MULTS_1_18(36)(PERCISION downto 1));
			MULTS_2_9(37)<=signed(MULTS_1_17(37)(PERCISION) & MULTS_1_17(37)(PERCISION downto 1))+signed(MULTS_1_18(37)(PERCISION) & MULTS_1_18(37)(PERCISION downto 1));
			MULTS_2_9(38)<=signed(MULTS_1_17(38)(PERCISION) & MULTS_1_17(38)(PERCISION downto 1))+signed(MULTS_1_18(38)(PERCISION) & MULTS_1_18(38)(PERCISION downto 1));
			MULTS_2_9(39)<=signed(MULTS_1_17(39)(PERCISION) & MULTS_1_17(39)(PERCISION downto 1))+signed(MULTS_1_18(39)(PERCISION) & MULTS_1_18(39)(PERCISION downto 1));
			MULTS_2_9(40)<=signed(MULTS_1_17(40)(PERCISION) & MULTS_1_17(40)(PERCISION downto 1))+signed(MULTS_1_18(40)(PERCISION) & MULTS_1_18(40)(PERCISION downto 1));
			MULTS_2_9(41)<=signed(MULTS_1_17(41)(PERCISION) & MULTS_1_17(41)(PERCISION downto 1))+signed(MULTS_1_18(41)(PERCISION) & MULTS_1_18(41)(PERCISION downto 1));
			MULTS_2_9(42)<=signed(MULTS_1_17(42)(PERCISION) & MULTS_1_17(42)(PERCISION downto 1))+signed(MULTS_1_18(42)(PERCISION) & MULTS_1_18(42)(PERCISION downto 1));
			MULTS_2_9(43)<=signed(MULTS_1_17(43)(PERCISION) & MULTS_1_17(43)(PERCISION downto 1))+signed(MULTS_1_18(43)(PERCISION) & MULTS_1_18(43)(PERCISION downto 1));
			MULTS_2_9(44)<=signed(MULTS_1_17(44)(PERCISION) & MULTS_1_17(44)(PERCISION downto 1))+signed(MULTS_1_18(44)(PERCISION) & MULTS_1_18(44)(PERCISION downto 1));
			MULTS_2_9(45)<=signed(MULTS_1_17(45)(PERCISION) & MULTS_1_17(45)(PERCISION downto 1))+signed(MULTS_1_18(45)(PERCISION) & MULTS_1_18(45)(PERCISION downto 1));
			MULTS_2_9(46)<=signed(MULTS_1_17(46)(PERCISION) & MULTS_1_17(46)(PERCISION downto 1))+signed(MULTS_1_18(46)(PERCISION) & MULTS_1_18(46)(PERCISION downto 1));
			MULTS_2_9(47)<=signed(MULTS_1_17(47)(PERCISION) & MULTS_1_17(47)(PERCISION downto 1))+signed(MULTS_1_18(47)(PERCISION) & MULTS_1_18(47)(PERCISION downto 1));
			MULTS_2_9(48)<=signed(MULTS_1_17(48)(PERCISION) & MULTS_1_17(48)(PERCISION downto 1))+signed(MULTS_1_18(48)(PERCISION) & MULTS_1_18(48)(PERCISION downto 1));
			MULTS_2_9(49)<=signed(MULTS_1_17(49)(PERCISION) & MULTS_1_17(49)(PERCISION downto 1))+signed(MULTS_1_18(49)(PERCISION) & MULTS_1_18(49)(PERCISION downto 1));
			MULTS_2_9(50)<=signed(MULTS_1_17(50)(PERCISION) & MULTS_1_17(50)(PERCISION downto 1))+signed(MULTS_1_18(50)(PERCISION) & MULTS_1_18(50)(PERCISION downto 1));
			MULTS_2_9(51)<=signed(MULTS_1_17(51)(PERCISION) & MULTS_1_17(51)(PERCISION downto 1))+signed(MULTS_1_18(51)(PERCISION) & MULTS_1_18(51)(PERCISION downto 1));
			MULTS_2_9(52)<=signed(MULTS_1_17(52)(PERCISION) & MULTS_1_17(52)(PERCISION downto 1))+signed(MULTS_1_18(52)(PERCISION) & MULTS_1_18(52)(PERCISION downto 1));
			MULTS_2_9(53)<=signed(MULTS_1_17(53)(PERCISION) & MULTS_1_17(53)(PERCISION downto 1))+signed(MULTS_1_18(53)(PERCISION) & MULTS_1_18(53)(PERCISION downto 1));
			MULTS_2_9(54)<=signed(MULTS_1_17(54)(PERCISION) & MULTS_1_17(54)(PERCISION downto 1))+signed(MULTS_1_18(54)(PERCISION) & MULTS_1_18(54)(PERCISION downto 1));
			MULTS_2_9(55)<=signed(MULTS_1_17(55)(PERCISION) & MULTS_1_17(55)(PERCISION downto 1))+signed(MULTS_1_18(55)(PERCISION) & MULTS_1_18(55)(PERCISION downto 1));
			MULTS_2_9(56)<=signed(MULTS_1_17(56)(PERCISION) & MULTS_1_17(56)(PERCISION downto 1))+signed(MULTS_1_18(56)(PERCISION) & MULTS_1_18(56)(PERCISION downto 1));
			MULTS_2_9(57)<=signed(MULTS_1_17(57)(PERCISION) & MULTS_1_17(57)(PERCISION downto 1))+signed(MULTS_1_18(57)(PERCISION) & MULTS_1_18(57)(PERCISION downto 1));
			MULTS_2_9(58)<=signed(MULTS_1_17(58)(PERCISION) & MULTS_1_17(58)(PERCISION downto 1))+signed(MULTS_1_18(58)(PERCISION) & MULTS_1_18(58)(PERCISION downto 1));
			MULTS_2_9(59)<=signed(MULTS_1_17(59)(PERCISION) & MULTS_1_17(59)(PERCISION downto 1))+signed(MULTS_1_18(59)(PERCISION) & MULTS_1_18(59)(PERCISION downto 1));
			MULTS_2_9(60)<=signed(MULTS_1_17(60)(PERCISION) & MULTS_1_17(60)(PERCISION downto 1))+signed(MULTS_1_18(60)(PERCISION) & MULTS_1_18(60)(PERCISION downto 1));
			MULTS_2_9(61)<=signed(MULTS_1_17(61)(PERCISION) & MULTS_1_17(61)(PERCISION downto 1))+signed(MULTS_1_18(61)(PERCISION) & MULTS_1_18(61)(PERCISION downto 1));
			MULTS_2_9(62)<=signed(MULTS_1_17(62)(PERCISION) & MULTS_1_17(62)(PERCISION downto 1))+signed(MULTS_1_18(62)(PERCISION) & MULTS_1_18(62)(PERCISION downto 1));
			MULTS_2_9(63)<=signed(MULTS_1_17(63)(PERCISION) & MULTS_1_17(63)(PERCISION downto 1))+signed(MULTS_1_18(63)(PERCISION) & MULTS_1_18(63)(PERCISION downto 1));
			MULTS_2_9(64)<=signed(MULTS_1_17(64)(PERCISION) & MULTS_1_17(64)(PERCISION downto 1))+signed(MULTS_1_18(64)(PERCISION) & MULTS_1_18(64)(PERCISION downto 1));
			MULTS_2_9(65)<=signed(MULTS_1_17(65)(PERCISION) & MULTS_1_17(65)(PERCISION downto 1))+signed(MULTS_1_18(65)(PERCISION) & MULTS_1_18(65)(PERCISION downto 1));
			MULTS_2_9(66)<=signed(MULTS_1_17(66)(PERCISION) & MULTS_1_17(66)(PERCISION downto 1))+signed(MULTS_1_18(66)(PERCISION) & MULTS_1_18(66)(PERCISION downto 1));
			MULTS_2_9(67)<=signed(MULTS_1_17(67)(PERCISION) & MULTS_1_17(67)(PERCISION downto 1))+signed(MULTS_1_18(67)(PERCISION) & MULTS_1_18(67)(PERCISION downto 1));
			MULTS_2_9(68)<=signed(MULTS_1_17(68)(PERCISION) & MULTS_1_17(68)(PERCISION downto 1))+signed(MULTS_1_18(68)(PERCISION) & MULTS_1_18(68)(PERCISION downto 1));
			MULTS_2_9(69)<=signed(MULTS_1_17(69)(PERCISION) & MULTS_1_17(69)(PERCISION downto 1))+signed(MULTS_1_18(69)(PERCISION) & MULTS_1_18(69)(PERCISION downto 1));
			MULTS_2_9(70)<=signed(MULTS_1_17(70)(PERCISION) & MULTS_1_17(70)(PERCISION downto 1))+signed(MULTS_1_18(70)(PERCISION) & MULTS_1_18(70)(PERCISION downto 1));
			MULTS_2_9(71)<=signed(MULTS_1_17(71)(PERCISION) & MULTS_1_17(71)(PERCISION downto 1))+signed(MULTS_1_18(71)(PERCISION) & MULTS_1_18(71)(PERCISION downto 1));
			MULTS_2_9(72)<=signed(MULTS_1_17(72)(PERCISION) & MULTS_1_17(72)(PERCISION downto 1))+signed(MULTS_1_18(72)(PERCISION) & MULTS_1_18(72)(PERCISION downto 1));
			MULTS_2_9(73)<=signed(MULTS_1_17(73)(PERCISION) & MULTS_1_17(73)(PERCISION downto 1))+signed(MULTS_1_18(73)(PERCISION) & MULTS_1_18(73)(PERCISION downto 1));
			MULTS_2_9(74)<=signed(MULTS_1_17(74)(PERCISION) & MULTS_1_17(74)(PERCISION downto 1))+signed(MULTS_1_18(74)(PERCISION) & MULTS_1_18(74)(PERCISION downto 1));
			MULTS_2_9(75)<=signed(MULTS_1_17(75)(PERCISION) & MULTS_1_17(75)(PERCISION downto 1))+signed(MULTS_1_18(75)(PERCISION) & MULTS_1_18(75)(PERCISION downto 1));
			MULTS_2_9(76)<=signed(MULTS_1_17(76)(PERCISION) & MULTS_1_17(76)(PERCISION downto 1))+signed(MULTS_1_18(76)(PERCISION) & MULTS_1_18(76)(PERCISION downto 1));
			MULTS_2_9(77)<=signed(MULTS_1_17(77)(PERCISION) & MULTS_1_17(77)(PERCISION downto 1))+signed(MULTS_1_18(77)(PERCISION) & MULTS_1_18(77)(PERCISION downto 1));
			MULTS_2_9(78)<=signed(MULTS_1_17(78)(PERCISION) & MULTS_1_17(78)(PERCISION downto 1))+signed(MULTS_1_18(78)(PERCISION) & MULTS_1_18(78)(PERCISION downto 1));
			MULTS_2_9(79)<=signed(MULTS_1_17(79)(PERCISION) & MULTS_1_17(79)(PERCISION downto 1))+signed(MULTS_1_18(79)(PERCISION) & MULTS_1_18(79)(PERCISION downto 1));
			MULTS_2_9(80)<=signed(MULTS_1_17(80)(PERCISION) & MULTS_1_17(80)(PERCISION downto 1))+signed(MULTS_1_18(80)(PERCISION) & MULTS_1_18(80)(PERCISION downto 1));
			MULTS_2_9(81)<=signed(MULTS_1_17(81)(PERCISION) & MULTS_1_17(81)(PERCISION downto 1))+signed(MULTS_1_18(81)(PERCISION) & MULTS_1_18(81)(PERCISION downto 1));
			MULTS_2_9(82)<=signed(MULTS_1_17(82)(PERCISION) & MULTS_1_17(82)(PERCISION downto 1))+signed(MULTS_1_18(82)(PERCISION) & MULTS_1_18(82)(PERCISION downto 1));
			MULTS_2_9(83)<=signed(MULTS_1_17(83)(PERCISION) & MULTS_1_17(83)(PERCISION downto 1))+signed(MULTS_1_18(83)(PERCISION) & MULTS_1_18(83)(PERCISION downto 1));

			MULTS_2_10(0)<=signed(MULTS_1_19(0)(PERCISION) & MULTS_1_19(0)(PERCISION downto 1))+signed(MULTS_1_20(0)(PERCISION) & MULTS_1_20(0)(PERCISION downto 1));
			MULTS_2_10(1)<=signed(MULTS_1_19(1)(PERCISION) & MULTS_1_19(1)(PERCISION downto 1))+signed(MULTS_1_20(1)(PERCISION) & MULTS_1_20(1)(PERCISION downto 1));
			MULTS_2_10(2)<=signed(MULTS_1_19(2)(PERCISION) & MULTS_1_19(2)(PERCISION downto 1))+signed(MULTS_1_20(2)(PERCISION) & MULTS_1_20(2)(PERCISION downto 1));
			MULTS_2_10(3)<=signed(MULTS_1_19(3)(PERCISION) & MULTS_1_19(3)(PERCISION downto 1))+signed(MULTS_1_20(3)(PERCISION) & MULTS_1_20(3)(PERCISION downto 1));
			MULTS_2_10(4)<=signed(MULTS_1_19(4)(PERCISION) & MULTS_1_19(4)(PERCISION downto 1))+signed(MULTS_1_20(4)(PERCISION) & MULTS_1_20(4)(PERCISION downto 1));
			MULTS_2_10(5)<=signed(MULTS_1_19(5)(PERCISION) & MULTS_1_19(5)(PERCISION downto 1))+signed(MULTS_1_20(5)(PERCISION) & MULTS_1_20(5)(PERCISION downto 1));
			MULTS_2_10(6)<=signed(MULTS_1_19(6)(PERCISION) & MULTS_1_19(6)(PERCISION downto 1))+signed(MULTS_1_20(6)(PERCISION) & MULTS_1_20(6)(PERCISION downto 1));
			MULTS_2_10(7)<=signed(MULTS_1_19(7)(PERCISION) & MULTS_1_19(7)(PERCISION downto 1))+signed(MULTS_1_20(7)(PERCISION) & MULTS_1_20(7)(PERCISION downto 1));
			MULTS_2_10(8)<=signed(MULTS_1_19(8)(PERCISION) & MULTS_1_19(8)(PERCISION downto 1))+signed(MULTS_1_20(8)(PERCISION) & MULTS_1_20(8)(PERCISION downto 1));
			MULTS_2_10(9)<=signed(MULTS_1_19(9)(PERCISION) & MULTS_1_19(9)(PERCISION downto 1))+signed(MULTS_1_20(9)(PERCISION) & MULTS_1_20(9)(PERCISION downto 1));
			MULTS_2_10(10)<=signed(MULTS_1_19(10)(PERCISION) & MULTS_1_19(10)(PERCISION downto 1))+signed(MULTS_1_20(10)(PERCISION) & MULTS_1_20(10)(PERCISION downto 1));
			MULTS_2_10(11)<=signed(MULTS_1_19(11)(PERCISION) & MULTS_1_19(11)(PERCISION downto 1))+signed(MULTS_1_20(11)(PERCISION) & MULTS_1_20(11)(PERCISION downto 1));
			MULTS_2_10(12)<=signed(MULTS_1_19(12)(PERCISION) & MULTS_1_19(12)(PERCISION downto 1))+signed(MULTS_1_20(12)(PERCISION) & MULTS_1_20(12)(PERCISION downto 1));
			MULTS_2_10(13)<=signed(MULTS_1_19(13)(PERCISION) & MULTS_1_19(13)(PERCISION downto 1))+signed(MULTS_1_20(13)(PERCISION) & MULTS_1_20(13)(PERCISION downto 1));
			MULTS_2_10(14)<=signed(MULTS_1_19(14)(PERCISION) & MULTS_1_19(14)(PERCISION downto 1))+signed(MULTS_1_20(14)(PERCISION) & MULTS_1_20(14)(PERCISION downto 1));
			MULTS_2_10(15)<=signed(MULTS_1_19(15)(PERCISION) & MULTS_1_19(15)(PERCISION downto 1))+signed(MULTS_1_20(15)(PERCISION) & MULTS_1_20(15)(PERCISION downto 1));
			MULTS_2_10(16)<=signed(MULTS_1_19(16)(PERCISION) & MULTS_1_19(16)(PERCISION downto 1))+signed(MULTS_1_20(16)(PERCISION) & MULTS_1_20(16)(PERCISION downto 1));
			MULTS_2_10(17)<=signed(MULTS_1_19(17)(PERCISION) & MULTS_1_19(17)(PERCISION downto 1))+signed(MULTS_1_20(17)(PERCISION) & MULTS_1_20(17)(PERCISION downto 1));
			MULTS_2_10(18)<=signed(MULTS_1_19(18)(PERCISION) & MULTS_1_19(18)(PERCISION downto 1))+signed(MULTS_1_20(18)(PERCISION) & MULTS_1_20(18)(PERCISION downto 1));
			MULTS_2_10(19)<=signed(MULTS_1_19(19)(PERCISION) & MULTS_1_19(19)(PERCISION downto 1))+signed(MULTS_1_20(19)(PERCISION) & MULTS_1_20(19)(PERCISION downto 1));
			MULTS_2_10(20)<=signed(MULTS_1_19(20)(PERCISION) & MULTS_1_19(20)(PERCISION downto 1))+signed(MULTS_1_20(20)(PERCISION) & MULTS_1_20(20)(PERCISION downto 1));
			MULTS_2_10(21)<=signed(MULTS_1_19(21)(PERCISION) & MULTS_1_19(21)(PERCISION downto 1))+signed(MULTS_1_20(21)(PERCISION) & MULTS_1_20(21)(PERCISION downto 1));
			MULTS_2_10(22)<=signed(MULTS_1_19(22)(PERCISION) & MULTS_1_19(22)(PERCISION downto 1))+signed(MULTS_1_20(22)(PERCISION) & MULTS_1_20(22)(PERCISION downto 1));
			MULTS_2_10(23)<=signed(MULTS_1_19(23)(PERCISION) & MULTS_1_19(23)(PERCISION downto 1))+signed(MULTS_1_20(23)(PERCISION) & MULTS_1_20(23)(PERCISION downto 1));
			MULTS_2_10(24)<=signed(MULTS_1_19(24)(PERCISION) & MULTS_1_19(24)(PERCISION downto 1))+signed(MULTS_1_20(24)(PERCISION) & MULTS_1_20(24)(PERCISION downto 1));
			MULTS_2_10(25)<=signed(MULTS_1_19(25)(PERCISION) & MULTS_1_19(25)(PERCISION downto 1))+signed(MULTS_1_20(25)(PERCISION) & MULTS_1_20(25)(PERCISION downto 1));
			MULTS_2_10(26)<=signed(MULTS_1_19(26)(PERCISION) & MULTS_1_19(26)(PERCISION downto 1))+signed(MULTS_1_20(26)(PERCISION) & MULTS_1_20(26)(PERCISION downto 1));
			MULTS_2_10(27)<=signed(MULTS_1_19(27)(PERCISION) & MULTS_1_19(27)(PERCISION downto 1))+signed(MULTS_1_20(27)(PERCISION) & MULTS_1_20(27)(PERCISION downto 1));
			MULTS_2_10(28)<=signed(MULTS_1_19(28)(PERCISION) & MULTS_1_19(28)(PERCISION downto 1))+signed(MULTS_1_20(28)(PERCISION) & MULTS_1_20(28)(PERCISION downto 1));
			MULTS_2_10(29)<=signed(MULTS_1_19(29)(PERCISION) & MULTS_1_19(29)(PERCISION downto 1))+signed(MULTS_1_20(29)(PERCISION) & MULTS_1_20(29)(PERCISION downto 1));
			MULTS_2_10(30)<=signed(MULTS_1_19(30)(PERCISION) & MULTS_1_19(30)(PERCISION downto 1))+signed(MULTS_1_20(30)(PERCISION) & MULTS_1_20(30)(PERCISION downto 1));
			MULTS_2_10(31)<=signed(MULTS_1_19(31)(PERCISION) & MULTS_1_19(31)(PERCISION downto 1))+signed(MULTS_1_20(31)(PERCISION) & MULTS_1_20(31)(PERCISION downto 1));
			MULTS_2_10(32)<=signed(MULTS_1_19(32)(PERCISION) & MULTS_1_19(32)(PERCISION downto 1))+signed(MULTS_1_20(32)(PERCISION) & MULTS_1_20(32)(PERCISION downto 1));
			MULTS_2_10(33)<=signed(MULTS_1_19(33)(PERCISION) & MULTS_1_19(33)(PERCISION downto 1))+signed(MULTS_1_20(33)(PERCISION) & MULTS_1_20(33)(PERCISION downto 1));
			MULTS_2_10(34)<=signed(MULTS_1_19(34)(PERCISION) & MULTS_1_19(34)(PERCISION downto 1))+signed(MULTS_1_20(34)(PERCISION) & MULTS_1_20(34)(PERCISION downto 1));
			MULTS_2_10(35)<=signed(MULTS_1_19(35)(PERCISION) & MULTS_1_19(35)(PERCISION downto 1))+signed(MULTS_1_20(35)(PERCISION) & MULTS_1_20(35)(PERCISION downto 1));
			MULTS_2_10(36)<=signed(MULTS_1_19(36)(PERCISION) & MULTS_1_19(36)(PERCISION downto 1))+signed(MULTS_1_20(36)(PERCISION) & MULTS_1_20(36)(PERCISION downto 1));
			MULTS_2_10(37)<=signed(MULTS_1_19(37)(PERCISION) & MULTS_1_19(37)(PERCISION downto 1))+signed(MULTS_1_20(37)(PERCISION) & MULTS_1_20(37)(PERCISION downto 1));
			MULTS_2_10(38)<=signed(MULTS_1_19(38)(PERCISION) & MULTS_1_19(38)(PERCISION downto 1))+signed(MULTS_1_20(38)(PERCISION) & MULTS_1_20(38)(PERCISION downto 1));
			MULTS_2_10(39)<=signed(MULTS_1_19(39)(PERCISION) & MULTS_1_19(39)(PERCISION downto 1))+signed(MULTS_1_20(39)(PERCISION) & MULTS_1_20(39)(PERCISION downto 1));
			MULTS_2_10(40)<=signed(MULTS_1_19(40)(PERCISION) & MULTS_1_19(40)(PERCISION downto 1))+signed(MULTS_1_20(40)(PERCISION) & MULTS_1_20(40)(PERCISION downto 1));
			MULTS_2_10(41)<=signed(MULTS_1_19(41)(PERCISION) & MULTS_1_19(41)(PERCISION downto 1))+signed(MULTS_1_20(41)(PERCISION) & MULTS_1_20(41)(PERCISION downto 1));
			MULTS_2_10(42)<=signed(MULTS_1_19(42)(PERCISION) & MULTS_1_19(42)(PERCISION downto 1))+signed(MULTS_1_20(42)(PERCISION) & MULTS_1_20(42)(PERCISION downto 1));
			MULTS_2_10(43)<=signed(MULTS_1_19(43)(PERCISION) & MULTS_1_19(43)(PERCISION downto 1))+signed(MULTS_1_20(43)(PERCISION) & MULTS_1_20(43)(PERCISION downto 1));
			MULTS_2_10(44)<=signed(MULTS_1_19(44)(PERCISION) & MULTS_1_19(44)(PERCISION downto 1))+signed(MULTS_1_20(44)(PERCISION) & MULTS_1_20(44)(PERCISION downto 1));
			MULTS_2_10(45)<=signed(MULTS_1_19(45)(PERCISION) & MULTS_1_19(45)(PERCISION downto 1))+signed(MULTS_1_20(45)(PERCISION) & MULTS_1_20(45)(PERCISION downto 1));
			MULTS_2_10(46)<=signed(MULTS_1_19(46)(PERCISION) & MULTS_1_19(46)(PERCISION downto 1))+signed(MULTS_1_20(46)(PERCISION) & MULTS_1_20(46)(PERCISION downto 1));
			MULTS_2_10(47)<=signed(MULTS_1_19(47)(PERCISION) & MULTS_1_19(47)(PERCISION downto 1))+signed(MULTS_1_20(47)(PERCISION) & MULTS_1_20(47)(PERCISION downto 1));
			MULTS_2_10(48)<=signed(MULTS_1_19(48)(PERCISION) & MULTS_1_19(48)(PERCISION downto 1))+signed(MULTS_1_20(48)(PERCISION) & MULTS_1_20(48)(PERCISION downto 1));
			MULTS_2_10(49)<=signed(MULTS_1_19(49)(PERCISION) & MULTS_1_19(49)(PERCISION downto 1))+signed(MULTS_1_20(49)(PERCISION) & MULTS_1_20(49)(PERCISION downto 1));
			MULTS_2_10(50)<=signed(MULTS_1_19(50)(PERCISION) & MULTS_1_19(50)(PERCISION downto 1))+signed(MULTS_1_20(50)(PERCISION) & MULTS_1_20(50)(PERCISION downto 1));
			MULTS_2_10(51)<=signed(MULTS_1_19(51)(PERCISION) & MULTS_1_19(51)(PERCISION downto 1))+signed(MULTS_1_20(51)(PERCISION) & MULTS_1_20(51)(PERCISION downto 1));
			MULTS_2_10(52)<=signed(MULTS_1_19(52)(PERCISION) & MULTS_1_19(52)(PERCISION downto 1))+signed(MULTS_1_20(52)(PERCISION) & MULTS_1_20(52)(PERCISION downto 1));
			MULTS_2_10(53)<=signed(MULTS_1_19(53)(PERCISION) & MULTS_1_19(53)(PERCISION downto 1))+signed(MULTS_1_20(53)(PERCISION) & MULTS_1_20(53)(PERCISION downto 1));
			MULTS_2_10(54)<=signed(MULTS_1_19(54)(PERCISION) & MULTS_1_19(54)(PERCISION downto 1))+signed(MULTS_1_20(54)(PERCISION) & MULTS_1_20(54)(PERCISION downto 1));
			MULTS_2_10(55)<=signed(MULTS_1_19(55)(PERCISION) & MULTS_1_19(55)(PERCISION downto 1))+signed(MULTS_1_20(55)(PERCISION) & MULTS_1_20(55)(PERCISION downto 1));
			MULTS_2_10(56)<=signed(MULTS_1_19(56)(PERCISION) & MULTS_1_19(56)(PERCISION downto 1))+signed(MULTS_1_20(56)(PERCISION) & MULTS_1_20(56)(PERCISION downto 1));
			MULTS_2_10(57)<=signed(MULTS_1_19(57)(PERCISION) & MULTS_1_19(57)(PERCISION downto 1))+signed(MULTS_1_20(57)(PERCISION) & MULTS_1_20(57)(PERCISION downto 1));
			MULTS_2_10(58)<=signed(MULTS_1_19(58)(PERCISION) & MULTS_1_19(58)(PERCISION downto 1))+signed(MULTS_1_20(58)(PERCISION) & MULTS_1_20(58)(PERCISION downto 1));
			MULTS_2_10(59)<=signed(MULTS_1_19(59)(PERCISION) & MULTS_1_19(59)(PERCISION downto 1))+signed(MULTS_1_20(59)(PERCISION) & MULTS_1_20(59)(PERCISION downto 1));
			MULTS_2_10(60)<=signed(MULTS_1_19(60)(PERCISION) & MULTS_1_19(60)(PERCISION downto 1))+signed(MULTS_1_20(60)(PERCISION) & MULTS_1_20(60)(PERCISION downto 1));
			MULTS_2_10(61)<=signed(MULTS_1_19(61)(PERCISION) & MULTS_1_19(61)(PERCISION downto 1))+signed(MULTS_1_20(61)(PERCISION) & MULTS_1_20(61)(PERCISION downto 1));
			MULTS_2_10(62)<=signed(MULTS_1_19(62)(PERCISION) & MULTS_1_19(62)(PERCISION downto 1))+signed(MULTS_1_20(62)(PERCISION) & MULTS_1_20(62)(PERCISION downto 1));
			MULTS_2_10(63)<=signed(MULTS_1_19(63)(PERCISION) & MULTS_1_19(63)(PERCISION downto 1))+signed(MULTS_1_20(63)(PERCISION) & MULTS_1_20(63)(PERCISION downto 1));
			MULTS_2_10(64)<=signed(MULTS_1_19(64)(PERCISION) & MULTS_1_19(64)(PERCISION downto 1))+signed(MULTS_1_20(64)(PERCISION) & MULTS_1_20(64)(PERCISION downto 1));
			MULTS_2_10(65)<=signed(MULTS_1_19(65)(PERCISION) & MULTS_1_19(65)(PERCISION downto 1))+signed(MULTS_1_20(65)(PERCISION) & MULTS_1_20(65)(PERCISION downto 1));
			MULTS_2_10(66)<=signed(MULTS_1_19(66)(PERCISION) & MULTS_1_19(66)(PERCISION downto 1))+signed(MULTS_1_20(66)(PERCISION) & MULTS_1_20(66)(PERCISION downto 1));
			MULTS_2_10(67)<=signed(MULTS_1_19(67)(PERCISION) & MULTS_1_19(67)(PERCISION downto 1))+signed(MULTS_1_20(67)(PERCISION) & MULTS_1_20(67)(PERCISION downto 1));
			MULTS_2_10(68)<=signed(MULTS_1_19(68)(PERCISION) & MULTS_1_19(68)(PERCISION downto 1))+signed(MULTS_1_20(68)(PERCISION) & MULTS_1_20(68)(PERCISION downto 1));
			MULTS_2_10(69)<=signed(MULTS_1_19(69)(PERCISION) & MULTS_1_19(69)(PERCISION downto 1))+signed(MULTS_1_20(69)(PERCISION) & MULTS_1_20(69)(PERCISION downto 1));
			MULTS_2_10(70)<=signed(MULTS_1_19(70)(PERCISION) & MULTS_1_19(70)(PERCISION downto 1))+signed(MULTS_1_20(70)(PERCISION) & MULTS_1_20(70)(PERCISION downto 1));
			MULTS_2_10(71)<=signed(MULTS_1_19(71)(PERCISION) & MULTS_1_19(71)(PERCISION downto 1))+signed(MULTS_1_20(71)(PERCISION) & MULTS_1_20(71)(PERCISION downto 1));
			MULTS_2_10(72)<=signed(MULTS_1_19(72)(PERCISION) & MULTS_1_19(72)(PERCISION downto 1))+signed(MULTS_1_20(72)(PERCISION) & MULTS_1_20(72)(PERCISION downto 1));
			MULTS_2_10(73)<=signed(MULTS_1_19(73)(PERCISION) & MULTS_1_19(73)(PERCISION downto 1))+signed(MULTS_1_20(73)(PERCISION) & MULTS_1_20(73)(PERCISION downto 1));
			MULTS_2_10(74)<=signed(MULTS_1_19(74)(PERCISION) & MULTS_1_19(74)(PERCISION downto 1))+signed(MULTS_1_20(74)(PERCISION) & MULTS_1_20(74)(PERCISION downto 1));
			MULTS_2_10(75)<=signed(MULTS_1_19(75)(PERCISION) & MULTS_1_19(75)(PERCISION downto 1))+signed(MULTS_1_20(75)(PERCISION) & MULTS_1_20(75)(PERCISION downto 1));
			MULTS_2_10(76)<=signed(MULTS_1_19(76)(PERCISION) & MULTS_1_19(76)(PERCISION downto 1))+signed(MULTS_1_20(76)(PERCISION) & MULTS_1_20(76)(PERCISION downto 1));
			MULTS_2_10(77)<=signed(MULTS_1_19(77)(PERCISION) & MULTS_1_19(77)(PERCISION downto 1))+signed(MULTS_1_20(77)(PERCISION) & MULTS_1_20(77)(PERCISION downto 1));
			MULTS_2_10(78)<=signed(MULTS_1_19(78)(PERCISION) & MULTS_1_19(78)(PERCISION downto 1))+signed(MULTS_1_20(78)(PERCISION) & MULTS_1_20(78)(PERCISION downto 1));
			MULTS_2_10(79)<=signed(MULTS_1_19(79)(PERCISION) & MULTS_1_19(79)(PERCISION downto 1))+signed(MULTS_1_20(79)(PERCISION) & MULTS_1_20(79)(PERCISION downto 1));
			MULTS_2_10(80)<=signed(MULTS_1_19(80)(PERCISION) & MULTS_1_19(80)(PERCISION downto 1))+signed(MULTS_1_20(80)(PERCISION) & MULTS_1_20(80)(PERCISION downto 1));
			MULTS_2_10(81)<=signed(MULTS_1_19(81)(PERCISION) & MULTS_1_19(81)(PERCISION downto 1))+signed(MULTS_1_20(81)(PERCISION) & MULTS_1_20(81)(PERCISION downto 1));
			MULTS_2_10(82)<=signed(MULTS_1_19(82)(PERCISION) & MULTS_1_19(82)(PERCISION downto 1))+signed(MULTS_1_20(82)(PERCISION) & MULTS_1_20(82)(PERCISION downto 1));
			MULTS_2_10(83)<=signed(MULTS_1_19(83)(PERCISION) & MULTS_1_19(83)(PERCISION downto 1))+signed(MULTS_1_20(83)(PERCISION) & MULTS_1_20(83)(PERCISION downto 1));

			MULTS_2_11(0)<=signed(MULTS_1_21(0)(PERCISION) & MULTS_1_21(0)(PERCISION downto 1))+signed(MULTS_1_22(0)(PERCISION) & MULTS_1_22(0)(PERCISION downto 1));
			MULTS_2_11(1)<=signed(MULTS_1_21(1)(PERCISION) & MULTS_1_21(1)(PERCISION downto 1))+signed(MULTS_1_22(1)(PERCISION) & MULTS_1_22(1)(PERCISION downto 1));
			MULTS_2_11(2)<=signed(MULTS_1_21(2)(PERCISION) & MULTS_1_21(2)(PERCISION downto 1))+signed(MULTS_1_22(2)(PERCISION) & MULTS_1_22(2)(PERCISION downto 1));
			MULTS_2_11(3)<=signed(MULTS_1_21(3)(PERCISION) & MULTS_1_21(3)(PERCISION downto 1))+signed(MULTS_1_22(3)(PERCISION) & MULTS_1_22(3)(PERCISION downto 1));
			MULTS_2_11(4)<=signed(MULTS_1_21(4)(PERCISION) & MULTS_1_21(4)(PERCISION downto 1))+signed(MULTS_1_22(4)(PERCISION) & MULTS_1_22(4)(PERCISION downto 1));
			MULTS_2_11(5)<=signed(MULTS_1_21(5)(PERCISION) & MULTS_1_21(5)(PERCISION downto 1))+signed(MULTS_1_22(5)(PERCISION) & MULTS_1_22(5)(PERCISION downto 1));
			MULTS_2_11(6)<=signed(MULTS_1_21(6)(PERCISION) & MULTS_1_21(6)(PERCISION downto 1))+signed(MULTS_1_22(6)(PERCISION) & MULTS_1_22(6)(PERCISION downto 1));
			MULTS_2_11(7)<=signed(MULTS_1_21(7)(PERCISION) & MULTS_1_21(7)(PERCISION downto 1))+signed(MULTS_1_22(7)(PERCISION) & MULTS_1_22(7)(PERCISION downto 1));
			MULTS_2_11(8)<=signed(MULTS_1_21(8)(PERCISION) & MULTS_1_21(8)(PERCISION downto 1))+signed(MULTS_1_22(8)(PERCISION) & MULTS_1_22(8)(PERCISION downto 1));
			MULTS_2_11(9)<=signed(MULTS_1_21(9)(PERCISION) & MULTS_1_21(9)(PERCISION downto 1))+signed(MULTS_1_22(9)(PERCISION) & MULTS_1_22(9)(PERCISION downto 1));
			MULTS_2_11(10)<=signed(MULTS_1_21(10)(PERCISION) & MULTS_1_21(10)(PERCISION downto 1))+signed(MULTS_1_22(10)(PERCISION) & MULTS_1_22(10)(PERCISION downto 1));
			MULTS_2_11(11)<=signed(MULTS_1_21(11)(PERCISION) & MULTS_1_21(11)(PERCISION downto 1))+signed(MULTS_1_22(11)(PERCISION) & MULTS_1_22(11)(PERCISION downto 1));
			MULTS_2_11(12)<=signed(MULTS_1_21(12)(PERCISION) & MULTS_1_21(12)(PERCISION downto 1))+signed(MULTS_1_22(12)(PERCISION) & MULTS_1_22(12)(PERCISION downto 1));
			MULTS_2_11(13)<=signed(MULTS_1_21(13)(PERCISION) & MULTS_1_21(13)(PERCISION downto 1))+signed(MULTS_1_22(13)(PERCISION) & MULTS_1_22(13)(PERCISION downto 1));
			MULTS_2_11(14)<=signed(MULTS_1_21(14)(PERCISION) & MULTS_1_21(14)(PERCISION downto 1))+signed(MULTS_1_22(14)(PERCISION) & MULTS_1_22(14)(PERCISION downto 1));
			MULTS_2_11(15)<=signed(MULTS_1_21(15)(PERCISION) & MULTS_1_21(15)(PERCISION downto 1))+signed(MULTS_1_22(15)(PERCISION) & MULTS_1_22(15)(PERCISION downto 1));
			MULTS_2_11(16)<=signed(MULTS_1_21(16)(PERCISION) & MULTS_1_21(16)(PERCISION downto 1))+signed(MULTS_1_22(16)(PERCISION) & MULTS_1_22(16)(PERCISION downto 1));
			MULTS_2_11(17)<=signed(MULTS_1_21(17)(PERCISION) & MULTS_1_21(17)(PERCISION downto 1))+signed(MULTS_1_22(17)(PERCISION) & MULTS_1_22(17)(PERCISION downto 1));
			MULTS_2_11(18)<=signed(MULTS_1_21(18)(PERCISION) & MULTS_1_21(18)(PERCISION downto 1))+signed(MULTS_1_22(18)(PERCISION) & MULTS_1_22(18)(PERCISION downto 1));
			MULTS_2_11(19)<=signed(MULTS_1_21(19)(PERCISION) & MULTS_1_21(19)(PERCISION downto 1))+signed(MULTS_1_22(19)(PERCISION) & MULTS_1_22(19)(PERCISION downto 1));
			MULTS_2_11(20)<=signed(MULTS_1_21(20)(PERCISION) & MULTS_1_21(20)(PERCISION downto 1))+signed(MULTS_1_22(20)(PERCISION) & MULTS_1_22(20)(PERCISION downto 1));
			MULTS_2_11(21)<=signed(MULTS_1_21(21)(PERCISION) & MULTS_1_21(21)(PERCISION downto 1))+signed(MULTS_1_22(21)(PERCISION) & MULTS_1_22(21)(PERCISION downto 1));
			MULTS_2_11(22)<=signed(MULTS_1_21(22)(PERCISION) & MULTS_1_21(22)(PERCISION downto 1))+signed(MULTS_1_22(22)(PERCISION) & MULTS_1_22(22)(PERCISION downto 1));
			MULTS_2_11(23)<=signed(MULTS_1_21(23)(PERCISION) & MULTS_1_21(23)(PERCISION downto 1))+signed(MULTS_1_22(23)(PERCISION) & MULTS_1_22(23)(PERCISION downto 1));
			MULTS_2_11(24)<=signed(MULTS_1_21(24)(PERCISION) & MULTS_1_21(24)(PERCISION downto 1))+signed(MULTS_1_22(24)(PERCISION) & MULTS_1_22(24)(PERCISION downto 1));
			MULTS_2_11(25)<=signed(MULTS_1_21(25)(PERCISION) & MULTS_1_21(25)(PERCISION downto 1))+signed(MULTS_1_22(25)(PERCISION) & MULTS_1_22(25)(PERCISION downto 1));
			MULTS_2_11(26)<=signed(MULTS_1_21(26)(PERCISION) & MULTS_1_21(26)(PERCISION downto 1))+signed(MULTS_1_22(26)(PERCISION) & MULTS_1_22(26)(PERCISION downto 1));
			MULTS_2_11(27)<=signed(MULTS_1_21(27)(PERCISION) & MULTS_1_21(27)(PERCISION downto 1))+signed(MULTS_1_22(27)(PERCISION) & MULTS_1_22(27)(PERCISION downto 1));
			MULTS_2_11(28)<=signed(MULTS_1_21(28)(PERCISION) & MULTS_1_21(28)(PERCISION downto 1))+signed(MULTS_1_22(28)(PERCISION) & MULTS_1_22(28)(PERCISION downto 1));
			MULTS_2_11(29)<=signed(MULTS_1_21(29)(PERCISION) & MULTS_1_21(29)(PERCISION downto 1))+signed(MULTS_1_22(29)(PERCISION) & MULTS_1_22(29)(PERCISION downto 1));
			MULTS_2_11(30)<=signed(MULTS_1_21(30)(PERCISION) & MULTS_1_21(30)(PERCISION downto 1))+signed(MULTS_1_22(30)(PERCISION) & MULTS_1_22(30)(PERCISION downto 1));
			MULTS_2_11(31)<=signed(MULTS_1_21(31)(PERCISION) & MULTS_1_21(31)(PERCISION downto 1))+signed(MULTS_1_22(31)(PERCISION) & MULTS_1_22(31)(PERCISION downto 1));
			MULTS_2_11(32)<=signed(MULTS_1_21(32)(PERCISION) & MULTS_1_21(32)(PERCISION downto 1))+signed(MULTS_1_22(32)(PERCISION) & MULTS_1_22(32)(PERCISION downto 1));
			MULTS_2_11(33)<=signed(MULTS_1_21(33)(PERCISION) & MULTS_1_21(33)(PERCISION downto 1))+signed(MULTS_1_22(33)(PERCISION) & MULTS_1_22(33)(PERCISION downto 1));
			MULTS_2_11(34)<=signed(MULTS_1_21(34)(PERCISION) & MULTS_1_21(34)(PERCISION downto 1))+signed(MULTS_1_22(34)(PERCISION) & MULTS_1_22(34)(PERCISION downto 1));
			MULTS_2_11(35)<=signed(MULTS_1_21(35)(PERCISION) & MULTS_1_21(35)(PERCISION downto 1))+signed(MULTS_1_22(35)(PERCISION) & MULTS_1_22(35)(PERCISION downto 1));
			MULTS_2_11(36)<=signed(MULTS_1_21(36)(PERCISION) & MULTS_1_21(36)(PERCISION downto 1))+signed(MULTS_1_22(36)(PERCISION) & MULTS_1_22(36)(PERCISION downto 1));
			MULTS_2_11(37)<=signed(MULTS_1_21(37)(PERCISION) & MULTS_1_21(37)(PERCISION downto 1))+signed(MULTS_1_22(37)(PERCISION) & MULTS_1_22(37)(PERCISION downto 1));
			MULTS_2_11(38)<=signed(MULTS_1_21(38)(PERCISION) & MULTS_1_21(38)(PERCISION downto 1))+signed(MULTS_1_22(38)(PERCISION) & MULTS_1_22(38)(PERCISION downto 1));
			MULTS_2_11(39)<=signed(MULTS_1_21(39)(PERCISION) & MULTS_1_21(39)(PERCISION downto 1))+signed(MULTS_1_22(39)(PERCISION) & MULTS_1_22(39)(PERCISION downto 1));
			MULTS_2_11(40)<=signed(MULTS_1_21(40)(PERCISION) & MULTS_1_21(40)(PERCISION downto 1))+signed(MULTS_1_22(40)(PERCISION) & MULTS_1_22(40)(PERCISION downto 1));
			MULTS_2_11(41)<=signed(MULTS_1_21(41)(PERCISION) & MULTS_1_21(41)(PERCISION downto 1))+signed(MULTS_1_22(41)(PERCISION) & MULTS_1_22(41)(PERCISION downto 1));
			MULTS_2_11(42)<=signed(MULTS_1_21(42)(PERCISION) & MULTS_1_21(42)(PERCISION downto 1))+signed(MULTS_1_22(42)(PERCISION) & MULTS_1_22(42)(PERCISION downto 1));
			MULTS_2_11(43)<=signed(MULTS_1_21(43)(PERCISION) & MULTS_1_21(43)(PERCISION downto 1))+signed(MULTS_1_22(43)(PERCISION) & MULTS_1_22(43)(PERCISION downto 1));
			MULTS_2_11(44)<=signed(MULTS_1_21(44)(PERCISION) & MULTS_1_21(44)(PERCISION downto 1))+signed(MULTS_1_22(44)(PERCISION) & MULTS_1_22(44)(PERCISION downto 1));
			MULTS_2_11(45)<=signed(MULTS_1_21(45)(PERCISION) & MULTS_1_21(45)(PERCISION downto 1))+signed(MULTS_1_22(45)(PERCISION) & MULTS_1_22(45)(PERCISION downto 1));
			MULTS_2_11(46)<=signed(MULTS_1_21(46)(PERCISION) & MULTS_1_21(46)(PERCISION downto 1))+signed(MULTS_1_22(46)(PERCISION) & MULTS_1_22(46)(PERCISION downto 1));
			MULTS_2_11(47)<=signed(MULTS_1_21(47)(PERCISION) & MULTS_1_21(47)(PERCISION downto 1))+signed(MULTS_1_22(47)(PERCISION) & MULTS_1_22(47)(PERCISION downto 1));
			MULTS_2_11(48)<=signed(MULTS_1_21(48)(PERCISION) & MULTS_1_21(48)(PERCISION downto 1))+signed(MULTS_1_22(48)(PERCISION) & MULTS_1_22(48)(PERCISION downto 1));
			MULTS_2_11(49)<=signed(MULTS_1_21(49)(PERCISION) & MULTS_1_21(49)(PERCISION downto 1))+signed(MULTS_1_22(49)(PERCISION) & MULTS_1_22(49)(PERCISION downto 1));
			MULTS_2_11(50)<=signed(MULTS_1_21(50)(PERCISION) & MULTS_1_21(50)(PERCISION downto 1))+signed(MULTS_1_22(50)(PERCISION) & MULTS_1_22(50)(PERCISION downto 1));
			MULTS_2_11(51)<=signed(MULTS_1_21(51)(PERCISION) & MULTS_1_21(51)(PERCISION downto 1))+signed(MULTS_1_22(51)(PERCISION) & MULTS_1_22(51)(PERCISION downto 1));
			MULTS_2_11(52)<=signed(MULTS_1_21(52)(PERCISION) & MULTS_1_21(52)(PERCISION downto 1))+signed(MULTS_1_22(52)(PERCISION) & MULTS_1_22(52)(PERCISION downto 1));
			MULTS_2_11(53)<=signed(MULTS_1_21(53)(PERCISION) & MULTS_1_21(53)(PERCISION downto 1))+signed(MULTS_1_22(53)(PERCISION) & MULTS_1_22(53)(PERCISION downto 1));
			MULTS_2_11(54)<=signed(MULTS_1_21(54)(PERCISION) & MULTS_1_21(54)(PERCISION downto 1))+signed(MULTS_1_22(54)(PERCISION) & MULTS_1_22(54)(PERCISION downto 1));
			MULTS_2_11(55)<=signed(MULTS_1_21(55)(PERCISION) & MULTS_1_21(55)(PERCISION downto 1))+signed(MULTS_1_22(55)(PERCISION) & MULTS_1_22(55)(PERCISION downto 1));
			MULTS_2_11(56)<=signed(MULTS_1_21(56)(PERCISION) & MULTS_1_21(56)(PERCISION downto 1))+signed(MULTS_1_22(56)(PERCISION) & MULTS_1_22(56)(PERCISION downto 1));
			MULTS_2_11(57)<=signed(MULTS_1_21(57)(PERCISION) & MULTS_1_21(57)(PERCISION downto 1))+signed(MULTS_1_22(57)(PERCISION) & MULTS_1_22(57)(PERCISION downto 1));
			MULTS_2_11(58)<=signed(MULTS_1_21(58)(PERCISION) & MULTS_1_21(58)(PERCISION downto 1))+signed(MULTS_1_22(58)(PERCISION) & MULTS_1_22(58)(PERCISION downto 1));
			MULTS_2_11(59)<=signed(MULTS_1_21(59)(PERCISION) & MULTS_1_21(59)(PERCISION downto 1))+signed(MULTS_1_22(59)(PERCISION) & MULTS_1_22(59)(PERCISION downto 1));
			MULTS_2_11(60)<=signed(MULTS_1_21(60)(PERCISION) & MULTS_1_21(60)(PERCISION downto 1))+signed(MULTS_1_22(60)(PERCISION) & MULTS_1_22(60)(PERCISION downto 1));
			MULTS_2_11(61)<=signed(MULTS_1_21(61)(PERCISION) & MULTS_1_21(61)(PERCISION downto 1))+signed(MULTS_1_22(61)(PERCISION) & MULTS_1_22(61)(PERCISION downto 1));
			MULTS_2_11(62)<=signed(MULTS_1_21(62)(PERCISION) & MULTS_1_21(62)(PERCISION downto 1))+signed(MULTS_1_22(62)(PERCISION) & MULTS_1_22(62)(PERCISION downto 1));
			MULTS_2_11(63)<=signed(MULTS_1_21(63)(PERCISION) & MULTS_1_21(63)(PERCISION downto 1))+signed(MULTS_1_22(63)(PERCISION) & MULTS_1_22(63)(PERCISION downto 1));
			MULTS_2_11(64)<=signed(MULTS_1_21(64)(PERCISION) & MULTS_1_21(64)(PERCISION downto 1))+signed(MULTS_1_22(64)(PERCISION) & MULTS_1_22(64)(PERCISION downto 1));
			MULTS_2_11(65)<=signed(MULTS_1_21(65)(PERCISION) & MULTS_1_21(65)(PERCISION downto 1))+signed(MULTS_1_22(65)(PERCISION) & MULTS_1_22(65)(PERCISION downto 1));
			MULTS_2_11(66)<=signed(MULTS_1_21(66)(PERCISION) & MULTS_1_21(66)(PERCISION downto 1))+signed(MULTS_1_22(66)(PERCISION) & MULTS_1_22(66)(PERCISION downto 1));
			MULTS_2_11(67)<=signed(MULTS_1_21(67)(PERCISION) & MULTS_1_21(67)(PERCISION downto 1))+signed(MULTS_1_22(67)(PERCISION) & MULTS_1_22(67)(PERCISION downto 1));
			MULTS_2_11(68)<=signed(MULTS_1_21(68)(PERCISION) & MULTS_1_21(68)(PERCISION downto 1))+signed(MULTS_1_22(68)(PERCISION) & MULTS_1_22(68)(PERCISION downto 1));
			MULTS_2_11(69)<=signed(MULTS_1_21(69)(PERCISION) & MULTS_1_21(69)(PERCISION downto 1))+signed(MULTS_1_22(69)(PERCISION) & MULTS_1_22(69)(PERCISION downto 1));
			MULTS_2_11(70)<=signed(MULTS_1_21(70)(PERCISION) & MULTS_1_21(70)(PERCISION downto 1))+signed(MULTS_1_22(70)(PERCISION) & MULTS_1_22(70)(PERCISION downto 1));
			MULTS_2_11(71)<=signed(MULTS_1_21(71)(PERCISION) & MULTS_1_21(71)(PERCISION downto 1))+signed(MULTS_1_22(71)(PERCISION) & MULTS_1_22(71)(PERCISION downto 1));
			MULTS_2_11(72)<=signed(MULTS_1_21(72)(PERCISION) & MULTS_1_21(72)(PERCISION downto 1))+signed(MULTS_1_22(72)(PERCISION) & MULTS_1_22(72)(PERCISION downto 1));
			MULTS_2_11(73)<=signed(MULTS_1_21(73)(PERCISION) & MULTS_1_21(73)(PERCISION downto 1))+signed(MULTS_1_22(73)(PERCISION) & MULTS_1_22(73)(PERCISION downto 1));
			MULTS_2_11(74)<=signed(MULTS_1_21(74)(PERCISION) & MULTS_1_21(74)(PERCISION downto 1))+signed(MULTS_1_22(74)(PERCISION) & MULTS_1_22(74)(PERCISION downto 1));
			MULTS_2_11(75)<=signed(MULTS_1_21(75)(PERCISION) & MULTS_1_21(75)(PERCISION downto 1))+signed(MULTS_1_22(75)(PERCISION) & MULTS_1_22(75)(PERCISION downto 1));
			MULTS_2_11(76)<=signed(MULTS_1_21(76)(PERCISION) & MULTS_1_21(76)(PERCISION downto 1))+signed(MULTS_1_22(76)(PERCISION) & MULTS_1_22(76)(PERCISION downto 1));
			MULTS_2_11(77)<=signed(MULTS_1_21(77)(PERCISION) & MULTS_1_21(77)(PERCISION downto 1))+signed(MULTS_1_22(77)(PERCISION) & MULTS_1_22(77)(PERCISION downto 1));
			MULTS_2_11(78)<=signed(MULTS_1_21(78)(PERCISION) & MULTS_1_21(78)(PERCISION downto 1))+signed(MULTS_1_22(78)(PERCISION) & MULTS_1_22(78)(PERCISION downto 1));
			MULTS_2_11(79)<=signed(MULTS_1_21(79)(PERCISION) & MULTS_1_21(79)(PERCISION downto 1))+signed(MULTS_1_22(79)(PERCISION) & MULTS_1_22(79)(PERCISION downto 1));
			MULTS_2_11(80)<=signed(MULTS_1_21(80)(PERCISION) & MULTS_1_21(80)(PERCISION downto 1))+signed(MULTS_1_22(80)(PERCISION) & MULTS_1_22(80)(PERCISION downto 1));
			MULTS_2_11(81)<=signed(MULTS_1_21(81)(PERCISION) & MULTS_1_21(81)(PERCISION downto 1))+signed(MULTS_1_22(81)(PERCISION) & MULTS_1_22(81)(PERCISION downto 1));
			MULTS_2_11(82)<=signed(MULTS_1_21(82)(PERCISION) & MULTS_1_21(82)(PERCISION downto 1))+signed(MULTS_1_22(82)(PERCISION) & MULTS_1_22(82)(PERCISION downto 1));
			MULTS_2_11(83)<=signed(MULTS_1_21(83)(PERCISION) & MULTS_1_21(83)(PERCISION downto 1))+signed(MULTS_1_22(83)(PERCISION) & MULTS_1_22(83)(PERCISION downto 1));

			MULTS_2_12(0)<=signed(MULTS_1_23(0)(PERCISION) & MULTS_1_23(0)(PERCISION downto 1))+signed(MULTS_1_24(0)(PERCISION) & MULTS_1_24(0)(PERCISION downto 1));
			MULTS_2_12(1)<=signed(MULTS_1_23(1)(PERCISION) & MULTS_1_23(1)(PERCISION downto 1))+signed(MULTS_1_24(1)(PERCISION) & MULTS_1_24(1)(PERCISION downto 1));
			MULTS_2_12(2)<=signed(MULTS_1_23(2)(PERCISION) & MULTS_1_23(2)(PERCISION downto 1))+signed(MULTS_1_24(2)(PERCISION) & MULTS_1_24(2)(PERCISION downto 1));
			MULTS_2_12(3)<=signed(MULTS_1_23(3)(PERCISION) & MULTS_1_23(3)(PERCISION downto 1))+signed(MULTS_1_24(3)(PERCISION) & MULTS_1_24(3)(PERCISION downto 1));
			MULTS_2_12(4)<=signed(MULTS_1_23(4)(PERCISION) & MULTS_1_23(4)(PERCISION downto 1))+signed(MULTS_1_24(4)(PERCISION) & MULTS_1_24(4)(PERCISION downto 1));
			MULTS_2_12(5)<=signed(MULTS_1_23(5)(PERCISION) & MULTS_1_23(5)(PERCISION downto 1))+signed(MULTS_1_24(5)(PERCISION) & MULTS_1_24(5)(PERCISION downto 1));
			MULTS_2_12(6)<=signed(MULTS_1_23(6)(PERCISION) & MULTS_1_23(6)(PERCISION downto 1))+signed(MULTS_1_24(6)(PERCISION) & MULTS_1_24(6)(PERCISION downto 1));
			MULTS_2_12(7)<=signed(MULTS_1_23(7)(PERCISION) & MULTS_1_23(7)(PERCISION downto 1))+signed(MULTS_1_24(7)(PERCISION) & MULTS_1_24(7)(PERCISION downto 1));
			MULTS_2_12(8)<=signed(MULTS_1_23(8)(PERCISION) & MULTS_1_23(8)(PERCISION downto 1))+signed(MULTS_1_24(8)(PERCISION) & MULTS_1_24(8)(PERCISION downto 1));
			MULTS_2_12(9)<=signed(MULTS_1_23(9)(PERCISION) & MULTS_1_23(9)(PERCISION downto 1))+signed(MULTS_1_24(9)(PERCISION) & MULTS_1_24(9)(PERCISION downto 1));
			MULTS_2_12(10)<=signed(MULTS_1_23(10)(PERCISION) & MULTS_1_23(10)(PERCISION downto 1))+signed(MULTS_1_24(10)(PERCISION) & MULTS_1_24(10)(PERCISION downto 1));
			MULTS_2_12(11)<=signed(MULTS_1_23(11)(PERCISION) & MULTS_1_23(11)(PERCISION downto 1))+signed(MULTS_1_24(11)(PERCISION) & MULTS_1_24(11)(PERCISION downto 1));
			MULTS_2_12(12)<=signed(MULTS_1_23(12)(PERCISION) & MULTS_1_23(12)(PERCISION downto 1))+signed(MULTS_1_24(12)(PERCISION) & MULTS_1_24(12)(PERCISION downto 1));
			MULTS_2_12(13)<=signed(MULTS_1_23(13)(PERCISION) & MULTS_1_23(13)(PERCISION downto 1))+signed(MULTS_1_24(13)(PERCISION) & MULTS_1_24(13)(PERCISION downto 1));
			MULTS_2_12(14)<=signed(MULTS_1_23(14)(PERCISION) & MULTS_1_23(14)(PERCISION downto 1))+signed(MULTS_1_24(14)(PERCISION) & MULTS_1_24(14)(PERCISION downto 1));
			MULTS_2_12(15)<=signed(MULTS_1_23(15)(PERCISION) & MULTS_1_23(15)(PERCISION downto 1))+signed(MULTS_1_24(15)(PERCISION) & MULTS_1_24(15)(PERCISION downto 1));
			MULTS_2_12(16)<=signed(MULTS_1_23(16)(PERCISION) & MULTS_1_23(16)(PERCISION downto 1))+signed(MULTS_1_24(16)(PERCISION) & MULTS_1_24(16)(PERCISION downto 1));
			MULTS_2_12(17)<=signed(MULTS_1_23(17)(PERCISION) & MULTS_1_23(17)(PERCISION downto 1))+signed(MULTS_1_24(17)(PERCISION) & MULTS_1_24(17)(PERCISION downto 1));
			MULTS_2_12(18)<=signed(MULTS_1_23(18)(PERCISION) & MULTS_1_23(18)(PERCISION downto 1))+signed(MULTS_1_24(18)(PERCISION) & MULTS_1_24(18)(PERCISION downto 1));
			MULTS_2_12(19)<=signed(MULTS_1_23(19)(PERCISION) & MULTS_1_23(19)(PERCISION downto 1))+signed(MULTS_1_24(19)(PERCISION) & MULTS_1_24(19)(PERCISION downto 1));
			MULTS_2_12(20)<=signed(MULTS_1_23(20)(PERCISION) & MULTS_1_23(20)(PERCISION downto 1))+signed(MULTS_1_24(20)(PERCISION) & MULTS_1_24(20)(PERCISION downto 1));
			MULTS_2_12(21)<=signed(MULTS_1_23(21)(PERCISION) & MULTS_1_23(21)(PERCISION downto 1))+signed(MULTS_1_24(21)(PERCISION) & MULTS_1_24(21)(PERCISION downto 1));
			MULTS_2_12(22)<=signed(MULTS_1_23(22)(PERCISION) & MULTS_1_23(22)(PERCISION downto 1))+signed(MULTS_1_24(22)(PERCISION) & MULTS_1_24(22)(PERCISION downto 1));
			MULTS_2_12(23)<=signed(MULTS_1_23(23)(PERCISION) & MULTS_1_23(23)(PERCISION downto 1))+signed(MULTS_1_24(23)(PERCISION) & MULTS_1_24(23)(PERCISION downto 1));
			MULTS_2_12(24)<=signed(MULTS_1_23(24)(PERCISION) & MULTS_1_23(24)(PERCISION downto 1))+signed(MULTS_1_24(24)(PERCISION) & MULTS_1_24(24)(PERCISION downto 1));
			MULTS_2_12(25)<=signed(MULTS_1_23(25)(PERCISION) & MULTS_1_23(25)(PERCISION downto 1))+signed(MULTS_1_24(25)(PERCISION) & MULTS_1_24(25)(PERCISION downto 1));
			MULTS_2_12(26)<=signed(MULTS_1_23(26)(PERCISION) & MULTS_1_23(26)(PERCISION downto 1))+signed(MULTS_1_24(26)(PERCISION) & MULTS_1_24(26)(PERCISION downto 1));
			MULTS_2_12(27)<=signed(MULTS_1_23(27)(PERCISION) & MULTS_1_23(27)(PERCISION downto 1))+signed(MULTS_1_24(27)(PERCISION) & MULTS_1_24(27)(PERCISION downto 1));
			MULTS_2_12(28)<=signed(MULTS_1_23(28)(PERCISION) & MULTS_1_23(28)(PERCISION downto 1))+signed(MULTS_1_24(28)(PERCISION) & MULTS_1_24(28)(PERCISION downto 1));
			MULTS_2_12(29)<=signed(MULTS_1_23(29)(PERCISION) & MULTS_1_23(29)(PERCISION downto 1))+signed(MULTS_1_24(29)(PERCISION) & MULTS_1_24(29)(PERCISION downto 1));
			MULTS_2_12(30)<=signed(MULTS_1_23(30)(PERCISION) & MULTS_1_23(30)(PERCISION downto 1))+signed(MULTS_1_24(30)(PERCISION) & MULTS_1_24(30)(PERCISION downto 1));
			MULTS_2_12(31)<=signed(MULTS_1_23(31)(PERCISION) & MULTS_1_23(31)(PERCISION downto 1))+signed(MULTS_1_24(31)(PERCISION) & MULTS_1_24(31)(PERCISION downto 1));
			MULTS_2_12(32)<=signed(MULTS_1_23(32)(PERCISION) & MULTS_1_23(32)(PERCISION downto 1))+signed(MULTS_1_24(32)(PERCISION) & MULTS_1_24(32)(PERCISION downto 1));
			MULTS_2_12(33)<=signed(MULTS_1_23(33)(PERCISION) & MULTS_1_23(33)(PERCISION downto 1))+signed(MULTS_1_24(33)(PERCISION) & MULTS_1_24(33)(PERCISION downto 1));
			MULTS_2_12(34)<=signed(MULTS_1_23(34)(PERCISION) & MULTS_1_23(34)(PERCISION downto 1))+signed(MULTS_1_24(34)(PERCISION) & MULTS_1_24(34)(PERCISION downto 1));
			MULTS_2_12(35)<=signed(MULTS_1_23(35)(PERCISION) & MULTS_1_23(35)(PERCISION downto 1))+signed(MULTS_1_24(35)(PERCISION) & MULTS_1_24(35)(PERCISION downto 1));
			MULTS_2_12(36)<=signed(MULTS_1_23(36)(PERCISION) & MULTS_1_23(36)(PERCISION downto 1))+signed(MULTS_1_24(36)(PERCISION) & MULTS_1_24(36)(PERCISION downto 1));
			MULTS_2_12(37)<=signed(MULTS_1_23(37)(PERCISION) & MULTS_1_23(37)(PERCISION downto 1))+signed(MULTS_1_24(37)(PERCISION) & MULTS_1_24(37)(PERCISION downto 1));
			MULTS_2_12(38)<=signed(MULTS_1_23(38)(PERCISION) & MULTS_1_23(38)(PERCISION downto 1))+signed(MULTS_1_24(38)(PERCISION) & MULTS_1_24(38)(PERCISION downto 1));
			MULTS_2_12(39)<=signed(MULTS_1_23(39)(PERCISION) & MULTS_1_23(39)(PERCISION downto 1))+signed(MULTS_1_24(39)(PERCISION) & MULTS_1_24(39)(PERCISION downto 1));
			MULTS_2_12(40)<=signed(MULTS_1_23(40)(PERCISION) & MULTS_1_23(40)(PERCISION downto 1))+signed(MULTS_1_24(40)(PERCISION) & MULTS_1_24(40)(PERCISION downto 1));
			MULTS_2_12(41)<=signed(MULTS_1_23(41)(PERCISION) & MULTS_1_23(41)(PERCISION downto 1))+signed(MULTS_1_24(41)(PERCISION) & MULTS_1_24(41)(PERCISION downto 1));
			MULTS_2_12(42)<=signed(MULTS_1_23(42)(PERCISION) & MULTS_1_23(42)(PERCISION downto 1))+signed(MULTS_1_24(42)(PERCISION) & MULTS_1_24(42)(PERCISION downto 1));
			MULTS_2_12(43)<=signed(MULTS_1_23(43)(PERCISION) & MULTS_1_23(43)(PERCISION downto 1))+signed(MULTS_1_24(43)(PERCISION) & MULTS_1_24(43)(PERCISION downto 1));
			MULTS_2_12(44)<=signed(MULTS_1_23(44)(PERCISION) & MULTS_1_23(44)(PERCISION downto 1))+signed(MULTS_1_24(44)(PERCISION) & MULTS_1_24(44)(PERCISION downto 1));
			MULTS_2_12(45)<=signed(MULTS_1_23(45)(PERCISION) & MULTS_1_23(45)(PERCISION downto 1))+signed(MULTS_1_24(45)(PERCISION) & MULTS_1_24(45)(PERCISION downto 1));
			MULTS_2_12(46)<=signed(MULTS_1_23(46)(PERCISION) & MULTS_1_23(46)(PERCISION downto 1))+signed(MULTS_1_24(46)(PERCISION) & MULTS_1_24(46)(PERCISION downto 1));
			MULTS_2_12(47)<=signed(MULTS_1_23(47)(PERCISION) & MULTS_1_23(47)(PERCISION downto 1))+signed(MULTS_1_24(47)(PERCISION) & MULTS_1_24(47)(PERCISION downto 1));
			MULTS_2_12(48)<=signed(MULTS_1_23(48)(PERCISION) & MULTS_1_23(48)(PERCISION downto 1))+signed(MULTS_1_24(48)(PERCISION) & MULTS_1_24(48)(PERCISION downto 1));
			MULTS_2_12(49)<=signed(MULTS_1_23(49)(PERCISION) & MULTS_1_23(49)(PERCISION downto 1))+signed(MULTS_1_24(49)(PERCISION) & MULTS_1_24(49)(PERCISION downto 1));
			MULTS_2_12(50)<=signed(MULTS_1_23(50)(PERCISION) & MULTS_1_23(50)(PERCISION downto 1))+signed(MULTS_1_24(50)(PERCISION) & MULTS_1_24(50)(PERCISION downto 1));
			MULTS_2_12(51)<=signed(MULTS_1_23(51)(PERCISION) & MULTS_1_23(51)(PERCISION downto 1))+signed(MULTS_1_24(51)(PERCISION) & MULTS_1_24(51)(PERCISION downto 1));
			MULTS_2_12(52)<=signed(MULTS_1_23(52)(PERCISION) & MULTS_1_23(52)(PERCISION downto 1))+signed(MULTS_1_24(52)(PERCISION) & MULTS_1_24(52)(PERCISION downto 1));
			MULTS_2_12(53)<=signed(MULTS_1_23(53)(PERCISION) & MULTS_1_23(53)(PERCISION downto 1))+signed(MULTS_1_24(53)(PERCISION) & MULTS_1_24(53)(PERCISION downto 1));
			MULTS_2_12(54)<=signed(MULTS_1_23(54)(PERCISION) & MULTS_1_23(54)(PERCISION downto 1))+signed(MULTS_1_24(54)(PERCISION) & MULTS_1_24(54)(PERCISION downto 1));
			MULTS_2_12(55)<=signed(MULTS_1_23(55)(PERCISION) & MULTS_1_23(55)(PERCISION downto 1))+signed(MULTS_1_24(55)(PERCISION) & MULTS_1_24(55)(PERCISION downto 1));
			MULTS_2_12(56)<=signed(MULTS_1_23(56)(PERCISION) & MULTS_1_23(56)(PERCISION downto 1))+signed(MULTS_1_24(56)(PERCISION) & MULTS_1_24(56)(PERCISION downto 1));
			MULTS_2_12(57)<=signed(MULTS_1_23(57)(PERCISION) & MULTS_1_23(57)(PERCISION downto 1))+signed(MULTS_1_24(57)(PERCISION) & MULTS_1_24(57)(PERCISION downto 1));
			MULTS_2_12(58)<=signed(MULTS_1_23(58)(PERCISION) & MULTS_1_23(58)(PERCISION downto 1))+signed(MULTS_1_24(58)(PERCISION) & MULTS_1_24(58)(PERCISION downto 1));
			MULTS_2_12(59)<=signed(MULTS_1_23(59)(PERCISION) & MULTS_1_23(59)(PERCISION downto 1))+signed(MULTS_1_24(59)(PERCISION) & MULTS_1_24(59)(PERCISION downto 1));
			MULTS_2_12(60)<=signed(MULTS_1_23(60)(PERCISION) & MULTS_1_23(60)(PERCISION downto 1))+signed(MULTS_1_24(60)(PERCISION) & MULTS_1_24(60)(PERCISION downto 1));
			MULTS_2_12(61)<=signed(MULTS_1_23(61)(PERCISION) & MULTS_1_23(61)(PERCISION downto 1))+signed(MULTS_1_24(61)(PERCISION) & MULTS_1_24(61)(PERCISION downto 1));
			MULTS_2_12(62)<=signed(MULTS_1_23(62)(PERCISION) & MULTS_1_23(62)(PERCISION downto 1))+signed(MULTS_1_24(62)(PERCISION) & MULTS_1_24(62)(PERCISION downto 1));
			MULTS_2_12(63)<=signed(MULTS_1_23(63)(PERCISION) & MULTS_1_23(63)(PERCISION downto 1))+signed(MULTS_1_24(63)(PERCISION) & MULTS_1_24(63)(PERCISION downto 1));
			MULTS_2_12(64)<=signed(MULTS_1_23(64)(PERCISION) & MULTS_1_23(64)(PERCISION downto 1))+signed(MULTS_1_24(64)(PERCISION) & MULTS_1_24(64)(PERCISION downto 1));
			MULTS_2_12(65)<=signed(MULTS_1_23(65)(PERCISION) & MULTS_1_23(65)(PERCISION downto 1))+signed(MULTS_1_24(65)(PERCISION) & MULTS_1_24(65)(PERCISION downto 1));
			MULTS_2_12(66)<=signed(MULTS_1_23(66)(PERCISION) & MULTS_1_23(66)(PERCISION downto 1))+signed(MULTS_1_24(66)(PERCISION) & MULTS_1_24(66)(PERCISION downto 1));
			MULTS_2_12(67)<=signed(MULTS_1_23(67)(PERCISION) & MULTS_1_23(67)(PERCISION downto 1))+signed(MULTS_1_24(67)(PERCISION) & MULTS_1_24(67)(PERCISION downto 1));
			MULTS_2_12(68)<=signed(MULTS_1_23(68)(PERCISION) & MULTS_1_23(68)(PERCISION downto 1))+signed(MULTS_1_24(68)(PERCISION) & MULTS_1_24(68)(PERCISION downto 1));
			MULTS_2_12(69)<=signed(MULTS_1_23(69)(PERCISION) & MULTS_1_23(69)(PERCISION downto 1))+signed(MULTS_1_24(69)(PERCISION) & MULTS_1_24(69)(PERCISION downto 1));
			MULTS_2_12(70)<=signed(MULTS_1_23(70)(PERCISION) & MULTS_1_23(70)(PERCISION downto 1))+signed(MULTS_1_24(70)(PERCISION) & MULTS_1_24(70)(PERCISION downto 1));
			MULTS_2_12(71)<=signed(MULTS_1_23(71)(PERCISION) & MULTS_1_23(71)(PERCISION downto 1))+signed(MULTS_1_24(71)(PERCISION) & MULTS_1_24(71)(PERCISION downto 1));
			MULTS_2_12(72)<=signed(MULTS_1_23(72)(PERCISION) & MULTS_1_23(72)(PERCISION downto 1))+signed(MULTS_1_24(72)(PERCISION) & MULTS_1_24(72)(PERCISION downto 1));
			MULTS_2_12(73)<=signed(MULTS_1_23(73)(PERCISION) & MULTS_1_23(73)(PERCISION downto 1))+signed(MULTS_1_24(73)(PERCISION) & MULTS_1_24(73)(PERCISION downto 1));
			MULTS_2_12(74)<=signed(MULTS_1_23(74)(PERCISION) & MULTS_1_23(74)(PERCISION downto 1))+signed(MULTS_1_24(74)(PERCISION) & MULTS_1_24(74)(PERCISION downto 1));
			MULTS_2_12(75)<=signed(MULTS_1_23(75)(PERCISION) & MULTS_1_23(75)(PERCISION downto 1))+signed(MULTS_1_24(75)(PERCISION) & MULTS_1_24(75)(PERCISION downto 1));
			MULTS_2_12(76)<=signed(MULTS_1_23(76)(PERCISION) & MULTS_1_23(76)(PERCISION downto 1))+signed(MULTS_1_24(76)(PERCISION) & MULTS_1_24(76)(PERCISION downto 1));
			MULTS_2_12(77)<=signed(MULTS_1_23(77)(PERCISION) & MULTS_1_23(77)(PERCISION downto 1))+signed(MULTS_1_24(77)(PERCISION) & MULTS_1_24(77)(PERCISION downto 1));
			MULTS_2_12(78)<=signed(MULTS_1_23(78)(PERCISION) & MULTS_1_23(78)(PERCISION downto 1))+signed(MULTS_1_24(78)(PERCISION) & MULTS_1_24(78)(PERCISION downto 1));
			MULTS_2_12(79)<=signed(MULTS_1_23(79)(PERCISION) & MULTS_1_23(79)(PERCISION downto 1))+signed(MULTS_1_24(79)(PERCISION) & MULTS_1_24(79)(PERCISION downto 1));
			MULTS_2_12(80)<=signed(MULTS_1_23(80)(PERCISION) & MULTS_1_23(80)(PERCISION downto 1))+signed(MULTS_1_24(80)(PERCISION) & MULTS_1_24(80)(PERCISION downto 1));
			MULTS_2_12(81)<=signed(MULTS_1_23(81)(PERCISION) & MULTS_1_23(81)(PERCISION downto 1))+signed(MULTS_1_24(81)(PERCISION) & MULTS_1_24(81)(PERCISION downto 1));
			MULTS_2_12(82)<=signed(MULTS_1_23(82)(PERCISION) & MULTS_1_23(82)(PERCISION downto 1))+signed(MULTS_1_24(82)(PERCISION) & MULTS_1_24(82)(PERCISION downto 1));
			MULTS_2_12(83)<=signed(MULTS_1_23(83)(PERCISION) & MULTS_1_23(83)(PERCISION downto 1))+signed(MULTS_1_24(83)(PERCISION) & MULTS_1_24(83)(PERCISION downto 1));

			MULTS_2_13(0)<=signed(MULTS_1_25(0)(PERCISION) & MULTS_1_25(0)(PERCISION downto 1))+signed(MULTS_1_26(0)(PERCISION) & MULTS_1_26(0)(PERCISION downto 1));
			MULTS_2_13(1)<=signed(MULTS_1_25(1)(PERCISION) & MULTS_1_25(1)(PERCISION downto 1))+signed(MULTS_1_26(1)(PERCISION) & MULTS_1_26(1)(PERCISION downto 1));
			MULTS_2_13(2)<=signed(MULTS_1_25(2)(PERCISION) & MULTS_1_25(2)(PERCISION downto 1))+signed(MULTS_1_26(2)(PERCISION) & MULTS_1_26(2)(PERCISION downto 1));
			MULTS_2_13(3)<=signed(MULTS_1_25(3)(PERCISION) & MULTS_1_25(3)(PERCISION downto 1))+signed(MULTS_1_26(3)(PERCISION) & MULTS_1_26(3)(PERCISION downto 1));
			MULTS_2_13(4)<=signed(MULTS_1_25(4)(PERCISION) & MULTS_1_25(4)(PERCISION downto 1))+signed(MULTS_1_26(4)(PERCISION) & MULTS_1_26(4)(PERCISION downto 1));
			MULTS_2_13(5)<=signed(MULTS_1_25(5)(PERCISION) & MULTS_1_25(5)(PERCISION downto 1))+signed(MULTS_1_26(5)(PERCISION) & MULTS_1_26(5)(PERCISION downto 1));
			MULTS_2_13(6)<=signed(MULTS_1_25(6)(PERCISION) & MULTS_1_25(6)(PERCISION downto 1))+signed(MULTS_1_26(6)(PERCISION) & MULTS_1_26(6)(PERCISION downto 1));
			MULTS_2_13(7)<=signed(MULTS_1_25(7)(PERCISION) & MULTS_1_25(7)(PERCISION downto 1))+signed(MULTS_1_26(7)(PERCISION) & MULTS_1_26(7)(PERCISION downto 1));
			MULTS_2_13(8)<=signed(MULTS_1_25(8)(PERCISION) & MULTS_1_25(8)(PERCISION downto 1))+signed(MULTS_1_26(8)(PERCISION) & MULTS_1_26(8)(PERCISION downto 1));
			MULTS_2_13(9)<=signed(MULTS_1_25(9)(PERCISION) & MULTS_1_25(9)(PERCISION downto 1))+signed(MULTS_1_26(9)(PERCISION) & MULTS_1_26(9)(PERCISION downto 1));
			MULTS_2_13(10)<=signed(MULTS_1_25(10)(PERCISION) & MULTS_1_25(10)(PERCISION downto 1))+signed(MULTS_1_26(10)(PERCISION) & MULTS_1_26(10)(PERCISION downto 1));
			MULTS_2_13(11)<=signed(MULTS_1_25(11)(PERCISION) & MULTS_1_25(11)(PERCISION downto 1))+signed(MULTS_1_26(11)(PERCISION) & MULTS_1_26(11)(PERCISION downto 1));
			MULTS_2_13(12)<=signed(MULTS_1_25(12)(PERCISION) & MULTS_1_25(12)(PERCISION downto 1))+signed(MULTS_1_26(12)(PERCISION) & MULTS_1_26(12)(PERCISION downto 1));
			MULTS_2_13(13)<=signed(MULTS_1_25(13)(PERCISION) & MULTS_1_25(13)(PERCISION downto 1))+signed(MULTS_1_26(13)(PERCISION) & MULTS_1_26(13)(PERCISION downto 1));
			MULTS_2_13(14)<=signed(MULTS_1_25(14)(PERCISION) & MULTS_1_25(14)(PERCISION downto 1))+signed(MULTS_1_26(14)(PERCISION) & MULTS_1_26(14)(PERCISION downto 1));
			MULTS_2_13(15)<=signed(MULTS_1_25(15)(PERCISION) & MULTS_1_25(15)(PERCISION downto 1))+signed(MULTS_1_26(15)(PERCISION) & MULTS_1_26(15)(PERCISION downto 1));
			MULTS_2_13(16)<=signed(MULTS_1_25(16)(PERCISION) & MULTS_1_25(16)(PERCISION downto 1))+signed(MULTS_1_26(16)(PERCISION) & MULTS_1_26(16)(PERCISION downto 1));
			MULTS_2_13(17)<=signed(MULTS_1_25(17)(PERCISION) & MULTS_1_25(17)(PERCISION downto 1))+signed(MULTS_1_26(17)(PERCISION) & MULTS_1_26(17)(PERCISION downto 1));
			MULTS_2_13(18)<=signed(MULTS_1_25(18)(PERCISION) & MULTS_1_25(18)(PERCISION downto 1))+signed(MULTS_1_26(18)(PERCISION) & MULTS_1_26(18)(PERCISION downto 1));
			MULTS_2_13(19)<=signed(MULTS_1_25(19)(PERCISION) & MULTS_1_25(19)(PERCISION downto 1))+signed(MULTS_1_26(19)(PERCISION) & MULTS_1_26(19)(PERCISION downto 1));
			MULTS_2_13(20)<=signed(MULTS_1_25(20)(PERCISION) & MULTS_1_25(20)(PERCISION downto 1))+signed(MULTS_1_26(20)(PERCISION) & MULTS_1_26(20)(PERCISION downto 1));
			MULTS_2_13(21)<=signed(MULTS_1_25(21)(PERCISION) & MULTS_1_25(21)(PERCISION downto 1))+signed(MULTS_1_26(21)(PERCISION) & MULTS_1_26(21)(PERCISION downto 1));
			MULTS_2_13(22)<=signed(MULTS_1_25(22)(PERCISION) & MULTS_1_25(22)(PERCISION downto 1))+signed(MULTS_1_26(22)(PERCISION) & MULTS_1_26(22)(PERCISION downto 1));
			MULTS_2_13(23)<=signed(MULTS_1_25(23)(PERCISION) & MULTS_1_25(23)(PERCISION downto 1))+signed(MULTS_1_26(23)(PERCISION) & MULTS_1_26(23)(PERCISION downto 1));
			MULTS_2_13(24)<=signed(MULTS_1_25(24)(PERCISION) & MULTS_1_25(24)(PERCISION downto 1))+signed(MULTS_1_26(24)(PERCISION) & MULTS_1_26(24)(PERCISION downto 1));
			MULTS_2_13(25)<=signed(MULTS_1_25(25)(PERCISION) & MULTS_1_25(25)(PERCISION downto 1))+signed(MULTS_1_26(25)(PERCISION) & MULTS_1_26(25)(PERCISION downto 1));
			MULTS_2_13(26)<=signed(MULTS_1_25(26)(PERCISION) & MULTS_1_25(26)(PERCISION downto 1))+signed(MULTS_1_26(26)(PERCISION) & MULTS_1_26(26)(PERCISION downto 1));
			MULTS_2_13(27)<=signed(MULTS_1_25(27)(PERCISION) & MULTS_1_25(27)(PERCISION downto 1))+signed(MULTS_1_26(27)(PERCISION) & MULTS_1_26(27)(PERCISION downto 1));
			MULTS_2_13(28)<=signed(MULTS_1_25(28)(PERCISION) & MULTS_1_25(28)(PERCISION downto 1))+signed(MULTS_1_26(28)(PERCISION) & MULTS_1_26(28)(PERCISION downto 1));
			MULTS_2_13(29)<=signed(MULTS_1_25(29)(PERCISION) & MULTS_1_25(29)(PERCISION downto 1))+signed(MULTS_1_26(29)(PERCISION) & MULTS_1_26(29)(PERCISION downto 1));
			MULTS_2_13(30)<=signed(MULTS_1_25(30)(PERCISION) & MULTS_1_25(30)(PERCISION downto 1))+signed(MULTS_1_26(30)(PERCISION) & MULTS_1_26(30)(PERCISION downto 1));
			MULTS_2_13(31)<=signed(MULTS_1_25(31)(PERCISION) & MULTS_1_25(31)(PERCISION downto 1))+signed(MULTS_1_26(31)(PERCISION) & MULTS_1_26(31)(PERCISION downto 1));
			MULTS_2_13(32)<=signed(MULTS_1_25(32)(PERCISION) & MULTS_1_25(32)(PERCISION downto 1))+signed(MULTS_1_26(32)(PERCISION) & MULTS_1_26(32)(PERCISION downto 1));
			MULTS_2_13(33)<=signed(MULTS_1_25(33)(PERCISION) & MULTS_1_25(33)(PERCISION downto 1))+signed(MULTS_1_26(33)(PERCISION) & MULTS_1_26(33)(PERCISION downto 1));
			MULTS_2_13(34)<=signed(MULTS_1_25(34)(PERCISION) & MULTS_1_25(34)(PERCISION downto 1))+signed(MULTS_1_26(34)(PERCISION) & MULTS_1_26(34)(PERCISION downto 1));
			MULTS_2_13(35)<=signed(MULTS_1_25(35)(PERCISION) & MULTS_1_25(35)(PERCISION downto 1))+signed(MULTS_1_26(35)(PERCISION) & MULTS_1_26(35)(PERCISION downto 1));
			MULTS_2_13(36)<=signed(MULTS_1_25(36)(PERCISION) & MULTS_1_25(36)(PERCISION downto 1))+signed(MULTS_1_26(36)(PERCISION) & MULTS_1_26(36)(PERCISION downto 1));
			MULTS_2_13(37)<=signed(MULTS_1_25(37)(PERCISION) & MULTS_1_25(37)(PERCISION downto 1))+signed(MULTS_1_26(37)(PERCISION) & MULTS_1_26(37)(PERCISION downto 1));
			MULTS_2_13(38)<=signed(MULTS_1_25(38)(PERCISION) & MULTS_1_25(38)(PERCISION downto 1))+signed(MULTS_1_26(38)(PERCISION) & MULTS_1_26(38)(PERCISION downto 1));
			MULTS_2_13(39)<=signed(MULTS_1_25(39)(PERCISION) & MULTS_1_25(39)(PERCISION downto 1))+signed(MULTS_1_26(39)(PERCISION) & MULTS_1_26(39)(PERCISION downto 1));
			MULTS_2_13(40)<=signed(MULTS_1_25(40)(PERCISION) & MULTS_1_25(40)(PERCISION downto 1))+signed(MULTS_1_26(40)(PERCISION) & MULTS_1_26(40)(PERCISION downto 1));
			MULTS_2_13(41)<=signed(MULTS_1_25(41)(PERCISION) & MULTS_1_25(41)(PERCISION downto 1))+signed(MULTS_1_26(41)(PERCISION) & MULTS_1_26(41)(PERCISION downto 1));
			MULTS_2_13(42)<=signed(MULTS_1_25(42)(PERCISION) & MULTS_1_25(42)(PERCISION downto 1))+signed(MULTS_1_26(42)(PERCISION) & MULTS_1_26(42)(PERCISION downto 1));
			MULTS_2_13(43)<=signed(MULTS_1_25(43)(PERCISION) & MULTS_1_25(43)(PERCISION downto 1))+signed(MULTS_1_26(43)(PERCISION) & MULTS_1_26(43)(PERCISION downto 1));
			MULTS_2_13(44)<=signed(MULTS_1_25(44)(PERCISION) & MULTS_1_25(44)(PERCISION downto 1))+signed(MULTS_1_26(44)(PERCISION) & MULTS_1_26(44)(PERCISION downto 1));
			MULTS_2_13(45)<=signed(MULTS_1_25(45)(PERCISION) & MULTS_1_25(45)(PERCISION downto 1))+signed(MULTS_1_26(45)(PERCISION) & MULTS_1_26(45)(PERCISION downto 1));
			MULTS_2_13(46)<=signed(MULTS_1_25(46)(PERCISION) & MULTS_1_25(46)(PERCISION downto 1))+signed(MULTS_1_26(46)(PERCISION) & MULTS_1_26(46)(PERCISION downto 1));
			MULTS_2_13(47)<=signed(MULTS_1_25(47)(PERCISION) & MULTS_1_25(47)(PERCISION downto 1))+signed(MULTS_1_26(47)(PERCISION) & MULTS_1_26(47)(PERCISION downto 1));
			MULTS_2_13(48)<=signed(MULTS_1_25(48)(PERCISION) & MULTS_1_25(48)(PERCISION downto 1))+signed(MULTS_1_26(48)(PERCISION) & MULTS_1_26(48)(PERCISION downto 1));
			MULTS_2_13(49)<=signed(MULTS_1_25(49)(PERCISION) & MULTS_1_25(49)(PERCISION downto 1))+signed(MULTS_1_26(49)(PERCISION) & MULTS_1_26(49)(PERCISION downto 1));
			MULTS_2_13(50)<=signed(MULTS_1_25(50)(PERCISION) & MULTS_1_25(50)(PERCISION downto 1))+signed(MULTS_1_26(50)(PERCISION) & MULTS_1_26(50)(PERCISION downto 1));
			MULTS_2_13(51)<=signed(MULTS_1_25(51)(PERCISION) & MULTS_1_25(51)(PERCISION downto 1))+signed(MULTS_1_26(51)(PERCISION) & MULTS_1_26(51)(PERCISION downto 1));
			MULTS_2_13(52)<=signed(MULTS_1_25(52)(PERCISION) & MULTS_1_25(52)(PERCISION downto 1))+signed(MULTS_1_26(52)(PERCISION) & MULTS_1_26(52)(PERCISION downto 1));
			MULTS_2_13(53)<=signed(MULTS_1_25(53)(PERCISION) & MULTS_1_25(53)(PERCISION downto 1))+signed(MULTS_1_26(53)(PERCISION) & MULTS_1_26(53)(PERCISION downto 1));
			MULTS_2_13(54)<=signed(MULTS_1_25(54)(PERCISION) & MULTS_1_25(54)(PERCISION downto 1))+signed(MULTS_1_26(54)(PERCISION) & MULTS_1_26(54)(PERCISION downto 1));
			MULTS_2_13(55)<=signed(MULTS_1_25(55)(PERCISION) & MULTS_1_25(55)(PERCISION downto 1))+signed(MULTS_1_26(55)(PERCISION) & MULTS_1_26(55)(PERCISION downto 1));
			MULTS_2_13(56)<=signed(MULTS_1_25(56)(PERCISION) & MULTS_1_25(56)(PERCISION downto 1))+signed(MULTS_1_26(56)(PERCISION) & MULTS_1_26(56)(PERCISION downto 1));
			MULTS_2_13(57)<=signed(MULTS_1_25(57)(PERCISION) & MULTS_1_25(57)(PERCISION downto 1))+signed(MULTS_1_26(57)(PERCISION) & MULTS_1_26(57)(PERCISION downto 1));
			MULTS_2_13(58)<=signed(MULTS_1_25(58)(PERCISION) & MULTS_1_25(58)(PERCISION downto 1))+signed(MULTS_1_26(58)(PERCISION) & MULTS_1_26(58)(PERCISION downto 1));
			MULTS_2_13(59)<=signed(MULTS_1_25(59)(PERCISION) & MULTS_1_25(59)(PERCISION downto 1))+signed(MULTS_1_26(59)(PERCISION) & MULTS_1_26(59)(PERCISION downto 1));
			MULTS_2_13(60)<=signed(MULTS_1_25(60)(PERCISION) & MULTS_1_25(60)(PERCISION downto 1))+signed(MULTS_1_26(60)(PERCISION) & MULTS_1_26(60)(PERCISION downto 1));
			MULTS_2_13(61)<=signed(MULTS_1_25(61)(PERCISION) & MULTS_1_25(61)(PERCISION downto 1))+signed(MULTS_1_26(61)(PERCISION) & MULTS_1_26(61)(PERCISION downto 1));
			MULTS_2_13(62)<=signed(MULTS_1_25(62)(PERCISION) & MULTS_1_25(62)(PERCISION downto 1))+signed(MULTS_1_26(62)(PERCISION) & MULTS_1_26(62)(PERCISION downto 1));
			MULTS_2_13(63)<=signed(MULTS_1_25(63)(PERCISION) & MULTS_1_25(63)(PERCISION downto 1))+signed(MULTS_1_26(63)(PERCISION) & MULTS_1_26(63)(PERCISION downto 1));
			MULTS_2_13(64)<=signed(MULTS_1_25(64)(PERCISION) & MULTS_1_25(64)(PERCISION downto 1))+signed(MULTS_1_26(64)(PERCISION) & MULTS_1_26(64)(PERCISION downto 1));
			MULTS_2_13(65)<=signed(MULTS_1_25(65)(PERCISION) & MULTS_1_25(65)(PERCISION downto 1))+signed(MULTS_1_26(65)(PERCISION) & MULTS_1_26(65)(PERCISION downto 1));
			MULTS_2_13(66)<=signed(MULTS_1_25(66)(PERCISION) & MULTS_1_25(66)(PERCISION downto 1))+signed(MULTS_1_26(66)(PERCISION) & MULTS_1_26(66)(PERCISION downto 1));
			MULTS_2_13(67)<=signed(MULTS_1_25(67)(PERCISION) & MULTS_1_25(67)(PERCISION downto 1))+signed(MULTS_1_26(67)(PERCISION) & MULTS_1_26(67)(PERCISION downto 1));
			MULTS_2_13(68)<=signed(MULTS_1_25(68)(PERCISION) & MULTS_1_25(68)(PERCISION downto 1))+signed(MULTS_1_26(68)(PERCISION) & MULTS_1_26(68)(PERCISION downto 1));
			MULTS_2_13(69)<=signed(MULTS_1_25(69)(PERCISION) & MULTS_1_25(69)(PERCISION downto 1))+signed(MULTS_1_26(69)(PERCISION) & MULTS_1_26(69)(PERCISION downto 1));
			MULTS_2_13(70)<=signed(MULTS_1_25(70)(PERCISION) & MULTS_1_25(70)(PERCISION downto 1))+signed(MULTS_1_26(70)(PERCISION) & MULTS_1_26(70)(PERCISION downto 1));
			MULTS_2_13(71)<=signed(MULTS_1_25(71)(PERCISION) & MULTS_1_25(71)(PERCISION downto 1))+signed(MULTS_1_26(71)(PERCISION) & MULTS_1_26(71)(PERCISION downto 1));
			MULTS_2_13(72)<=signed(MULTS_1_25(72)(PERCISION) & MULTS_1_25(72)(PERCISION downto 1))+signed(MULTS_1_26(72)(PERCISION) & MULTS_1_26(72)(PERCISION downto 1));
			MULTS_2_13(73)<=signed(MULTS_1_25(73)(PERCISION) & MULTS_1_25(73)(PERCISION downto 1))+signed(MULTS_1_26(73)(PERCISION) & MULTS_1_26(73)(PERCISION downto 1));
			MULTS_2_13(74)<=signed(MULTS_1_25(74)(PERCISION) & MULTS_1_25(74)(PERCISION downto 1))+signed(MULTS_1_26(74)(PERCISION) & MULTS_1_26(74)(PERCISION downto 1));
			MULTS_2_13(75)<=signed(MULTS_1_25(75)(PERCISION) & MULTS_1_25(75)(PERCISION downto 1))+signed(MULTS_1_26(75)(PERCISION) & MULTS_1_26(75)(PERCISION downto 1));
			MULTS_2_13(76)<=signed(MULTS_1_25(76)(PERCISION) & MULTS_1_25(76)(PERCISION downto 1))+signed(MULTS_1_26(76)(PERCISION) & MULTS_1_26(76)(PERCISION downto 1));
			MULTS_2_13(77)<=signed(MULTS_1_25(77)(PERCISION) & MULTS_1_25(77)(PERCISION downto 1))+signed(MULTS_1_26(77)(PERCISION) & MULTS_1_26(77)(PERCISION downto 1));
			MULTS_2_13(78)<=signed(MULTS_1_25(78)(PERCISION) & MULTS_1_25(78)(PERCISION downto 1))+signed(MULTS_1_26(78)(PERCISION) & MULTS_1_26(78)(PERCISION downto 1));
			MULTS_2_13(79)<=signed(MULTS_1_25(79)(PERCISION) & MULTS_1_25(79)(PERCISION downto 1))+signed(MULTS_1_26(79)(PERCISION) & MULTS_1_26(79)(PERCISION downto 1));
			MULTS_2_13(80)<=signed(MULTS_1_25(80)(PERCISION) & MULTS_1_25(80)(PERCISION downto 1))+signed(MULTS_1_26(80)(PERCISION) & MULTS_1_26(80)(PERCISION downto 1));
			MULTS_2_13(81)<=signed(MULTS_1_25(81)(PERCISION) & MULTS_1_25(81)(PERCISION downto 1))+signed(MULTS_1_26(81)(PERCISION) & MULTS_1_26(81)(PERCISION downto 1));
			MULTS_2_13(82)<=signed(MULTS_1_25(82)(PERCISION) & MULTS_1_25(82)(PERCISION downto 1))+signed(MULTS_1_26(82)(PERCISION) & MULTS_1_26(82)(PERCISION downto 1));
			MULTS_2_13(83)<=signed(MULTS_1_25(83)(PERCISION) & MULTS_1_25(83)(PERCISION downto 1))+signed(MULTS_1_26(83)(PERCISION) & MULTS_1_26(83)(PERCISION downto 1));

			MULTS_2_14(0)<=signed(MULTS_1_27(0)(PERCISION) & MULTS_1_27(0)(PERCISION downto 1))+signed(MULTS_1_28(0)(PERCISION) & MULTS_1_28(0)(PERCISION downto 1));
			MULTS_2_14(1)<=signed(MULTS_1_27(1)(PERCISION) & MULTS_1_27(1)(PERCISION downto 1))+signed(MULTS_1_28(1)(PERCISION) & MULTS_1_28(1)(PERCISION downto 1));
			MULTS_2_14(2)<=signed(MULTS_1_27(2)(PERCISION) & MULTS_1_27(2)(PERCISION downto 1))+signed(MULTS_1_28(2)(PERCISION) & MULTS_1_28(2)(PERCISION downto 1));
			MULTS_2_14(3)<=signed(MULTS_1_27(3)(PERCISION) & MULTS_1_27(3)(PERCISION downto 1))+signed(MULTS_1_28(3)(PERCISION) & MULTS_1_28(3)(PERCISION downto 1));
			MULTS_2_14(4)<=signed(MULTS_1_27(4)(PERCISION) & MULTS_1_27(4)(PERCISION downto 1))+signed(MULTS_1_28(4)(PERCISION) & MULTS_1_28(4)(PERCISION downto 1));
			MULTS_2_14(5)<=signed(MULTS_1_27(5)(PERCISION) & MULTS_1_27(5)(PERCISION downto 1))+signed(MULTS_1_28(5)(PERCISION) & MULTS_1_28(5)(PERCISION downto 1));
			MULTS_2_14(6)<=signed(MULTS_1_27(6)(PERCISION) & MULTS_1_27(6)(PERCISION downto 1))+signed(MULTS_1_28(6)(PERCISION) & MULTS_1_28(6)(PERCISION downto 1));
			MULTS_2_14(7)<=signed(MULTS_1_27(7)(PERCISION) & MULTS_1_27(7)(PERCISION downto 1))+signed(MULTS_1_28(7)(PERCISION) & MULTS_1_28(7)(PERCISION downto 1));
			MULTS_2_14(8)<=signed(MULTS_1_27(8)(PERCISION) & MULTS_1_27(8)(PERCISION downto 1))+signed(MULTS_1_28(8)(PERCISION) & MULTS_1_28(8)(PERCISION downto 1));
			MULTS_2_14(9)<=signed(MULTS_1_27(9)(PERCISION) & MULTS_1_27(9)(PERCISION downto 1))+signed(MULTS_1_28(9)(PERCISION) & MULTS_1_28(9)(PERCISION downto 1));
			MULTS_2_14(10)<=signed(MULTS_1_27(10)(PERCISION) & MULTS_1_27(10)(PERCISION downto 1))+signed(MULTS_1_28(10)(PERCISION) & MULTS_1_28(10)(PERCISION downto 1));
			MULTS_2_14(11)<=signed(MULTS_1_27(11)(PERCISION) & MULTS_1_27(11)(PERCISION downto 1))+signed(MULTS_1_28(11)(PERCISION) & MULTS_1_28(11)(PERCISION downto 1));
			MULTS_2_14(12)<=signed(MULTS_1_27(12)(PERCISION) & MULTS_1_27(12)(PERCISION downto 1))+signed(MULTS_1_28(12)(PERCISION) & MULTS_1_28(12)(PERCISION downto 1));
			MULTS_2_14(13)<=signed(MULTS_1_27(13)(PERCISION) & MULTS_1_27(13)(PERCISION downto 1))+signed(MULTS_1_28(13)(PERCISION) & MULTS_1_28(13)(PERCISION downto 1));
			MULTS_2_14(14)<=signed(MULTS_1_27(14)(PERCISION) & MULTS_1_27(14)(PERCISION downto 1))+signed(MULTS_1_28(14)(PERCISION) & MULTS_1_28(14)(PERCISION downto 1));
			MULTS_2_14(15)<=signed(MULTS_1_27(15)(PERCISION) & MULTS_1_27(15)(PERCISION downto 1))+signed(MULTS_1_28(15)(PERCISION) & MULTS_1_28(15)(PERCISION downto 1));
			MULTS_2_14(16)<=signed(MULTS_1_27(16)(PERCISION) & MULTS_1_27(16)(PERCISION downto 1))+signed(MULTS_1_28(16)(PERCISION) & MULTS_1_28(16)(PERCISION downto 1));
			MULTS_2_14(17)<=signed(MULTS_1_27(17)(PERCISION) & MULTS_1_27(17)(PERCISION downto 1))+signed(MULTS_1_28(17)(PERCISION) & MULTS_1_28(17)(PERCISION downto 1));
			MULTS_2_14(18)<=signed(MULTS_1_27(18)(PERCISION) & MULTS_1_27(18)(PERCISION downto 1))+signed(MULTS_1_28(18)(PERCISION) & MULTS_1_28(18)(PERCISION downto 1));
			MULTS_2_14(19)<=signed(MULTS_1_27(19)(PERCISION) & MULTS_1_27(19)(PERCISION downto 1))+signed(MULTS_1_28(19)(PERCISION) & MULTS_1_28(19)(PERCISION downto 1));
			MULTS_2_14(20)<=signed(MULTS_1_27(20)(PERCISION) & MULTS_1_27(20)(PERCISION downto 1))+signed(MULTS_1_28(20)(PERCISION) & MULTS_1_28(20)(PERCISION downto 1));
			MULTS_2_14(21)<=signed(MULTS_1_27(21)(PERCISION) & MULTS_1_27(21)(PERCISION downto 1))+signed(MULTS_1_28(21)(PERCISION) & MULTS_1_28(21)(PERCISION downto 1));
			MULTS_2_14(22)<=signed(MULTS_1_27(22)(PERCISION) & MULTS_1_27(22)(PERCISION downto 1))+signed(MULTS_1_28(22)(PERCISION) & MULTS_1_28(22)(PERCISION downto 1));
			MULTS_2_14(23)<=signed(MULTS_1_27(23)(PERCISION) & MULTS_1_27(23)(PERCISION downto 1))+signed(MULTS_1_28(23)(PERCISION) & MULTS_1_28(23)(PERCISION downto 1));
			MULTS_2_14(24)<=signed(MULTS_1_27(24)(PERCISION) & MULTS_1_27(24)(PERCISION downto 1))+signed(MULTS_1_28(24)(PERCISION) & MULTS_1_28(24)(PERCISION downto 1));
			MULTS_2_14(25)<=signed(MULTS_1_27(25)(PERCISION) & MULTS_1_27(25)(PERCISION downto 1))+signed(MULTS_1_28(25)(PERCISION) & MULTS_1_28(25)(PERCISION downto 1));
			MULTS_2_14(26)<=signed(MULTS_1_27(26)(PERCISION) & MULTS_1_27(26)(PERCISION downto 1))+signed(MULTS_1_28(26)(PERCISION) & MULTS_1_28(26)(PERCISION downto 1));
			MULTS_2_14(27)<=signed(MULTS_1_27(27)(PERCISION) & MULTS_1_27(27)(PERCISION downto 1))+signed(MULTS_1_28(27)(PERCISION) & MULTS_1_28(27)(PERCISION downto 1));
			MULTS_2_14(28)<=signed(MULTS_1_27(28)(PERCISION) & MULTS_1_27(28)(PERCISION downto 1))+signed(MULTS_1_28(28)(PERCISION) & MULTS_1_28(28)(PERCISION downto 1));
			MULTS_2_14(29)<=signed(MULTS_1_27(29)(PERCISION) & MULTS_1_27(29)(PERCISION downto 1))+signed(MULTS_1_28(29)(PERCISION) & MULTS_1_28(29)(PERCISION downto 1));
			MULTS_2_14(30)<=signed(MULTS_1_27(30)(PERCISION) & MULTS_1_27(30)(PERCISION downto 1))+signed(MULTS_1_28(30)(PERCISION) & MULTS_1_28(30)(PERCISION downto 1));
			MULTS_2_14(31)<=signed(MULTS_1_27(31)(PERCISION) & MULTS_1_27(31)(PERCISION downto 1))+signed(MULTS_1_28(31)(PERCISION) & MULTS_1_28(31)(PERCISION downto 1));
			MULTS_2_14(32)<=signed(MULTS_1_27(32)(PERCISION) & MULTS_1_27(32)(PERCISION downto 1))+signed(MULTS_1_28(32)(PERCISION) & MULTS_1_28(32)(PERCISION downto 1));
			MULTS_2_14(33)<=signed(MULTS_1_27(33)(PERCISION) & MULTS_1_27(33)(PERCISION downto 1))+signed(MULTS_1_28(33)(PERCISION) & MULTS_1_28(33)(PERCISION downto 1));
			MULTS_2_14(34)<=signed(MULTS_1_27(34)(PERCISION) & MULTS_1_27(34)(PERCISION downto 1))+signed(MULTS_1_28(34)(PERCISION) & MULTS_1_28(34)(PERCISION downto 1));
			MULTS_2_14(35)<=signed(MULTS_1_27(35)(PERCISION) & MULTS_1_27(35)(PERCISION downto 1))+signed(MULTS_1_28(35)(PERCISION) & MULTS_1_28(35)(PERCISION downto 1));
			MULTS_2_14(36)<=signed(MULTS_1_27(36)(PERCISION) & MULTS_1_27(36)(PERCISION downto 1))+signed(MULTS_1_28(36)(PERCISION) & MULTS_1_28(36)(PERCISION downto 1));
			MULTS_2_14(37)<=signed(MULTS_1_27(37)(PERCISION) & MULTS_1_27(37)(PERCISION downto 1))+signed(MULTS_1_28(37)(PERCISION) & MULTS_1_28(37)(PERCISION downto 1));
			MULTS_2_14(38)<=signed(MULTS_1_27(38)(PERCISION) & MULTS_1_27(38)(PERCISION downto 1))+signed(MULTS_1_28(38)(PERCISION) & MULTS_1_28(38)(PERCISION downto 1));
			MULTS_2_14(39)<=signed(MULTS_1_27(39)(PERCISION) & MULTS_1_27(39)(PERCISION downto 1))+signed(MULTS_1_28(39)(PERCISION) & MULTS_1_28(39)(PERCISION downto 1));
			MULTS_2_14(40)<=signed(MULTS_1_27(40)(PERCISION) & MULTS_1_27(40)(PERCISION downto 1))+signed(MULTS_1_28(40)(PERCISION) & MULTS_1_28(40)(PERCISION downto 1));
			MULTS_2_14(41)<=signed(MULTS_1_27(41)(PERCISION) & MULTS_1_27(41)(PERCISION downto 1))+signed(MULTS_1_28(41)(PERCISION) & MULTS_1_28(41)(PERCISION downto 1));
			MULTS_2_14(42)<=signed(MULTS_1_27(42)(PERCISION) & MULTS_1_27(42)(PERCISION downto 1))+signed(MULTS_1_28(42)(PERCISION) & MULTS_1_28(42)(PERCISION downto 1));
			MULTS_2_14(43)<=signed(MULTS_1_27(43)(PERCISION) & MULTS_1_27(43)(PERCISION downto 1))+signed(MULTS_1_28(43)(PERCISION) & MULTS_1_28(43)(PERCISION downto 1));
			MULTS_2_14(44)<=signed(MULTS_1_27(44)(PERCISION) & MULTS_1_27(44)(PERCISION downto 1))+signed(MULTS_1_28(44)(PERCISION) & MULTS_1_28(44)(PERCISION downto 1));
			MULTS_2_14(45)<=signed(MULTS_1_27(45)(PERCISION) & MULTS_1_27(45)(PERCISION downto 1))+signed(MULTS_1_28(45)(PERCISION) & MULTS_1_28(45)(PERCISION downto 1));
			MULTS_2_14(46)<=signed(MULTS_1_27(46)(PERCISION) & MULTS_1_27(46)(PERCISION downto 1))+signed(MULTS_1_28(46)(PERCISION) & MULTS_1_28(46)(PERCISION downto 1));
			MULTS_2_14(47)<=signed(MULTS_1_27(47)(PERCISION) & MULTS_1_27(47)(PERCISION downto 1))+signed(MULTS_1_28(47)(PERCISION) & MULTS_1_28(47)(PERCISION downto 1));
			MULTS_2_14(48)<=signed(MULTS_1_27(48)(PERCISION) & MULTS_1_27(48)(PERCISION downto 1))+signed(MULTS_1_28(48)(PERCISION) & MULTS_1_28(48)(PERCISION downto 1));
			MULTS_2_14(49)<=signed(MULTS_1_27(49)(PERCISION) & MULTS_1_27(49)(PERCISION downto 1))+signed(MULTS_1_28(49)(PERCISION) & MULTS_1_28(49)(PERCISION downto 1));
			MULTS_2_14(50)<=signed(MULTS_1_27(50)(PERCISION) & MULTS_1_27(50)(PERCISION downto 1))+signed(MULTS_1_28(50)(PERCISION) & MULTS_1_28(50)(PERCISION downto 1));
			MULTS_2_14(51)<=signed(MULTS_1_27(51)(PERCISION) & MULTS_1_27(51)(PERCISION downto 1))+signed(MULTS_1_28(51)(PERCISION) & MULTS_1_28(51)(PERCISION downto 1));
			MULTS_2_14(52)<=signed(MULTS_1_27(52)(PERCISION) & MULTS_1_27(52)(PERCISION downto 1))+signed(MULTS_1_28(52)(PERCISION) & MULTS_1_28(52)(PERCISION downto 1));
			MULTS_2_14(53)<=signed(MULTS_1_27(53)(PERCISION) & MULTS_1_27(53)(PERCISION downto 1))+signed(MULTS_1_28(53)(PERCISION) & MULTS_1_28(53)(PERCISION downto 1));
			MULTS_2_14(54)<=signed(MULTS_1_27(54)(PERCISION) & MULTS_1_27(54)(PERCISION downto 1))+signed(MULTS_1_28(54)(PERCISION) & MULTS_1_28(54)(PERCISION downto 1));
			MULTS_2_14(55)<=signed(MULTS_1_27(55)(PERCISION) & MULTS_1_27(55)(PERCISION downto 1))+signed(MULTS_1_28(55)(PERCISION) & MULTS_1_28(55)(PERCISION downto 1));
			MULTS_2_14(56)<=signed(MULTS_1_27(56)(PERCISION) & MULTS_1_27(56)(PERCISION downto 1))+signed(MULTS_1_28(56)(PERCISION) & MULTS_1_28(56)(PERCISION downto 1));
			MULTS_2_14(57)<=signed(MULTS_1_27(57)(PERCISION) & MULTS_1_27(57)(PERCISION downto 1))+signed(MULTS_1_28(57)(PERCISION) & MULTS_1_28(57)(PERCISION downto 1));
			MULTS_2_14(58)<=signed(MULTS_1_27(58)(PERCISION) & MULTS_1_27(58)(PERCISION downto 1))+signed(MULTS_1_28(58)(PERCISION) & MULTS_1_28(58)(PERCISION downto 1));
			MULTS_2_14(59)<=signed(MULTS_1_27(59)(PERCISION) & MULTS_1_27(59)(PERCISION downto 1))+signed(MULTS_1_28(59)(PERCISION) & MULTS_1_28(59)(PERCISION downto 1));
			MULTS_2_14(60)<=signed(MULTS_1_27(60)(PERCISION) & MULTS_1_27(60)(PERCISION downto 1))+signed(MULTS_1_28(60)(PERCISION) & MULTS_1_28(60)(PERCISION downto 1));
			MULTS_2_14(61)<=signed(MULTS_1_27(61)(PERCISION) & MULTS_1_27(61)(PERCISION downto 1))+signed(MULTS_1_28(61)(PERCISION) & MULTS_1_28(61)(PERCISION downto 1));
			MULTS_2_14(62)<=signed(MULTS_1_27(62)(PERCISION) & MULTS_1_27(62)(PERCISION downto 1))+signed(MULTS_1_28(62)(PERCISION) & MULTS_1_28(62)(PERCISION downto 1));
			MULTS_2_14(63)<=signed(MULTS_1_27(63)(PERCISION) & MULTS_1_27(63)(PERCISION downto 1))+signed(MULTS_1_28(63)(PERCISION) & MULTS_1_28(63)(PERCISION downto 1));
			MULTS_2_14(64)<=signed(MULTS_1_27(64)(PERCISION) & MULTS_1_27(64)(PERCISION downto 1))+signed(MULTS_1_28(64)(PERCISION) & MULTS_1_28(64)(PERCISION downto 1));
			MULTS_2_14(65)<=signed(MULTS_1_27(65)(PERCISION) & MULTS_1_27(65)(PERCISION downto 1))+signed(MULTS_1_28(65)(PERCISION) & MULTS_1_28(65)(PERCISION downto 1));
			MULTS_2_14(66)<=signed(MULTS_1_27(66)(PERCISION) & MULTS_1_27(66)(PERCISION downto 1))+signed(MULTS_1_28(66)(PERCISION) & MULTS_1_28(66)(PERCISION downto 1));
			MULTS_2_14(67)<=signed(MULTS_1_27(67)(PERCISION) & MULTS_1_27(67)(PERCISION downto 1))+signed(MULTS_1_28(67)(PERCISION) & MULTS_1_28(67)(PERCISION downto 1));
			MULTS_2_14(68)<=signed(MULTS_1_27(68)(PERCISION) & MULTS_1_27(68)(PERCISION downto 1))+signed(MULTS_1_28(68)(PERCISION) & MULTS_1_28(68)(PERCISION downto 1));
			MULTS_2_14(69)<=signed(MULTS_1_27(69)(PERCISION) & MULTS_1_27(69)(PERCISION downto 1))+signed(MULTS_1_28(69)(PERCISION) & MULTS_1_28(69)(PERCISION downto 1));
			MULTS_2_14(70)<=signed(MULTS_1_27(70)(PERCISION) & MULTS_1_27(70)(PERCISION downto 1))+signed(MULTS_1_28(70)(PERCISION) & MULTS_1_28(70)(PERCISION downto 1));
			MULTS_2_14(71)<=signed(MULTS_1_27(71)(PERCISION) & MULTS_1_27(71)(PERCISION downto 1))+signed(MULTS_1_28(71)(PERCISION) & MULTS_1_28(71)(PERCISION downto 1));
			MULTS_2_14(72)<=signed(MULTS_1_27(72)(PERCISION) & MULTS_1_27(72)(PERCISION downto 1))+signed(MULTS_1_28(72)(PERCISION) & MULTS_1_28(72)(PERCISION downto 1));
			MULTS_2_14(73)<=signed(MULTS_1_27(73)(PERCISION) & MULTS_1_27(73)(PERCISION downto 1))+signed(MULTS_1_28(73)(PERCISION) & MULTS_1_28(73)(PERCISION downto 1));
			MULTS_2_14(74)<=signed(MULTS_1_27(74)(PERCISION) & MULTS_1_27(74)(PERCISION downto 1))+signed(MULTS_1_28(74)(PERCISION) & MULTS_1_28(74)(PERCISION downto 1));
			MULTS_2_14(75)<=signed(MULTS_1_27(75)(PERCISION) & MULTS_1_27(75)(PERCISION downto 1))+signed(MULTS_1_28(75)(PERCISION) & MULTS_1_28(75)(PERCISION downto 1));
			MULTS_2_14(76)<=signed(MULTS_1_27(76)(PERCISION) & MULTS_1_27(76)(PERCISION downto 1))+signed(MULTS_1_28(76)(PERCISION) & MULTS_1_28(76)(PERCISION downto 1));
			MULTS_2_14(77)<=signed(MULTS_1_27(77)(PERCISION) & MULTS_1_27(77)(PERCISION downto 1))+signed(MULTS_1_28(77)(PERCISION) & MULTS_1_28(77)(PERCISION downto 1));
			MULTS_2_14(78)<=signed(MULTS_1_27(78)(PERCISION) & MULTS_1_27(78)(PERCISION downto 1))+signed(MULTS_1_28(78)(PERCISION) & MULTS_1_28(78)(PERCISION downto 1));
			MULTS_2_14(79)<=signed(MULTS_1_27(79)(PERCISION) & MULTS_1_27(79)(PERCISION downto 1))+signed(MULTS_1_28(79)(PERCISION) & MULTS_1_28(79)(PERCISION downto 1));
			MULTS_2_14(80)<=signed(MULTS_1_27(80)(PERCISION) & MULTS_1_27(80)(PERCISION downto 1))+signed(MULTS_1_28(80)(PERCISION) & MULTS_1_28(80)(PERCISION downto 1));
			MULTS_2_14(81)<=signed(MULTS_1_27(81)(PERCISION) & MULTS_1_27(81)(PERCISION downto 1))+signed(MULTS_1_28(81)(PERCISION) & MULTS_1_28(81)(PERCISION downto 1));
			MULTS_2_14(82)<=signed(MULTS_1_27(82)(PERCISION) & MULTS_1_27(82)(PERCISION downto 1))+signed(MULTS_1_28(82)(PERCISION) & MULTS_1_28(82)(PERCISION downto 1));
			MULTS_2_14(83)<=signed(MULTS_1_27(83)(PERCISION) & MULTS_1_27(83)(PERCISION downto 1))+signed(MULTS_1_28(83)(PERCISION) & MULTS_1_28(83)(PERCISION downto 1));

			MULTS_2_15(0)<=signed(MULTS_1_29(0)(PERCISION) & MULTS_1_29(0)(PERCISION downto 1))+signed(MULTS_1_30(0)(PERCISION) & MULTS_1_30(0)(PERCISION downto 1));
			MULTS_2_15(1)<=signed(MULTS_1_29(1)(PERCISION) & MULTS_1_29(1)(PERCISION downto 1))+signed(MULTS_1_30(1)(PERCISION) & MULTS_1_30(1)(PERCISION downto 1));
			MULTS_2_15(2)<=signed(MULTS_1_29(2)(PERCISION) & MULTS_1_29(2)(PERCISION downto 1))+signed(MULTS_1_30(2)(PERCISION) & MULTS_1_30(2)(PERCISION downto 1));
			MULTS_2_15(3)<=signed(MULTS_1_29(3)(PERCISION) & MULTS_1_29(3)(PERCISION downto 1))+signed(MULTS_1_30(3)(PERCISION) & MULTS_1_30(3)(PERCISION downto 1));
			MULTS_2_15(4)<=signed(MULTS_1_29(4)(PERCISION) & MULTS_1_29(4)(PERCISION downto 1))+signed(MULTS_1_30(4)(PERCISION) & MULTS_1_30(4)(PERCISION downto 1));
			MULTS_2_15(5)<=signed(MULTS_1_29(5)(PERCISION) & MULTS_1_29(5)(PERCISION downto 1))+signed(MULTS_1_30(5)(PERCISION) & MULTS_1_30(5)(PERCISION downto 1));
			MULTS_2_15(6)<=signed(MULTS_1_29(6)(PERCISION) & MULTS_1_29(6)(PERCISION downto 1))+signed(MULTS_1_30(6)(PERCISION) & MULTS_1_30(6)(PERCISION downto 1));
			MULTS_2_15(7)<=signed(MULTS_1_29(7)(PERCISION) & MULTS_1_29(7)(PERCISION downto 1))+signed(MULTS_1_30(7)(PERCISION) & MULTS_1_30(7)(PERCISION downto 1));
			MULTS_2_15(8)<=signed(MULTS_1_29(8)(PERCISION) & MULTS_1_29(8)(PERCISION downto 1))+signed(MULTS_1_30(8)(PERCISION) & MULTS_1_30(8)(PERCISION downto 1));
			MULTS_2_15(9)<=signed(MULTS_1_29(9)(PERCISION) & MULTS_1_29(9)(PERCISION downto 1))+signed(MULTS_1_30(9)(PERCISION) & MULTS_1_30(9)(PERCISION downto 1));
			MULTS_2_15(10)<=signed(MULTS_1_29(10)(PERCISION) & MULTS_1_29(10)(PERCISION downto 1))+signed(MULTS_1_30(10)(PERCISION) & MULTS_1_30(10)(PERCISION downto 1));
			MULTS_2_15(11)<=signed(MULTS_1_29(11)(PERCISION) & MULTS_1_29(11)(PERCISION downto 1))+signed(MULTS_1_30(11)(PERCISION) & MULTS_1_30(11)(PERCISION downto 1));
			MULTS_2_15(12)<=signed(MULTS_1_29(12)(PERCISION) & MULTS_1_29(12)(PERCISION downto 1))+signed(MULTS_1_30(12)(PERCISION) & MULTS_1_30(12)(PERCISION downto 1));
			MULTS_2_15(13)<=signed(MULTS_1_29(13)(PERCISION) & MULTS_1_29(13)(PERCISION downto 1))+signed(MULTS_1_30(13)(PERCISION) & MULTS_1_30(13)(PERCISION downto 1));
			MULTS_2_15(14)<=signed(MULTS_1_29(14)(PERCISION) & MULTS_1_29(14)(PERCISION downto 1))+signed(MULTS_1_30(14)(PERCISION) & MULTS_1_30(14)(PERCISION downto 1));
			MULTS_2_15(15)<=signed(MULTS_1_29(15)(PERCISION) & MULTS_1_29(15)(PERCISION downto 1))+signed(MULTS_1_30(15)(PERCISION) & MULTS_1_30(15)(PERCISION downto 1));
			MULTS_2_15(16)<=signed(MULTS_1_29(16)(PERCISION) & MULTS_1_29(16)(PERCISION downto 1))+signed(MULTS_1_30(16)(PERCISION) & MULTS_1_30(16)(PERCISION downto 1));
			MULTS_2_15(17)<=signed(MULTS_1_29(17)(PERCISION) & MULTS_1_29(17)(PERCISION downto 1))+signed(MULTS_1_30(17)(PERCISION) & MULTS_1_30(17)(PERCISION downto 1));
			MULTS_2_15(18)<=signed(MULTS_1_29(18)(PERCISION) & MULTS_1_29(18)(PERCISION downto 1))+signed(MULTS_1_30(18)(PERCISION) & MULTS_1_30(18)(PERCISION downto 1));
			MULTS_2_15(19)<=signed(MULTS_1_29(19)(PERCISION) & MULTS_1_29(19)(PERCISION downto 1))+signed(MULTS_1_30(19)(PERCISION) & MULTS_1_30(19)(PERCISION downto 1));
			MULTS_2_15(20)<=signed(MULTS_1_29(20)(PERCISION) & MULTS_1_29(20)(PERCISION downto 1))+signed(MULTS_1_30(20)(PERCISION) & MULTS_1_30(20)(PERCISION downto 1));
			MULTS_2_15(21)<=signed(MULTS_1_29(21)(PERCISION) & MULTS_1_29(21)(PERCISION downto 1))+signed(MULTS_1_30(21)(PERCISION) & MULTS_1_30(21)(PERCISION downto 1));
			MULTS_2_15(22)<=signed(MULTS_1_29(22)(PERCISION) & MULTS_1_29(22)(PERCISION downto 1))+signed(MULTS_1_30(22)(PERCISION) & MULTS_1_30(22)(PERCISION downto 1));
			MULTS_2_15(23)<=signed(MULTS_1_29(23)(PERCISION) & MULTS_1_29(23)(PERCISION downto 1))+signed(MULTS_1_30(23)(PERCISION) & MULTS_1_30(23)(PERCISION downto 1));
			MULTS_2_15(24)<=signed(MULTS_1_29(24)(PERCISION) & MULTS_1_29(24)(PERCISION downto 1))+signed(MULTS_1_30(24)(PERCISION) & MULTS_1_30(24)(PERCISION downto 1));
			MULTS_2_15(25)<=signed(MULTS_1_29(25)(PERCISION) & MULTS_1_29(25)(PERCISION downto 1))+signed(MULTS_1_30(25)(PERCISION) & MULTS_1_30(25)(PERCISION downto 1));
			MULTS_2_15(26)<=signed(MULTS_1_29(26)(PERCISION) & MULTS_1_29(26)(PERCISION downto 1))+signed(MULTS_1_30(26)(PERCISION) & MULTS_1_30(26)(PERCISION downto 1));
			MULTS_2_15(27)<=signed(MULTS_1_29(27)(PERCISION) & MULTS_1_29(27)(PERCISION downto 1))+signed(MULTS_1_30(27)(PERCISION) & MULTS_1_30(27)(PERCISION downto 1));
			MULTS_2_15(28)<=signed(MULTS_1_29(28)(PERCISION) & MULTS_1_29(28)(PERCISION downto 1))+signed(MULTS_1_30(28)(PERCISION) & MULTS_1_30(28)(PERCISION downto 1));
			MULTS_2_15(29)<=signed(MULTS_1_29(29)(PERCISION) & MULTS_1_29(29)(PERCISION downto 1))+signed(MULTS_1_30(29)(PERCISION) & MULTS_1_30(29)(PERCISION downto 1));
			MULTS_2_15(30)<=signed(MULTS_1_29(30)(PERCISION) & MULTS_1_29(30)(PERCISION downto 1))+signed(MULTS_1_30(30)(PERCISION) & MULTS_1_30(30)(PERCISION downto 1));
			MULTS_2_15(31)<=signed(MULTS_1_29(31)(PERCISION) & MULTS_1_29(31)(PERCISION downto 1))+signed(MULTS_1_30(31)(PERCISION) & MULTS_1_30(31)(PERCISION downto 1));
			MULTS_2_15(32)<=signed(MULTS_1_29(32)(PERCISION) & MULTS_1_29(32)(PERCISION downto 1))+signed(MULTS_1_30(32)(PERCISION) & MULTS_1_30(32)(PERCISION downto 1));
			MULTS_2_15(33)<=signed(MULTS_1_29(33)(PERCISION) & MULTS_1_29(33)(PERCISION downto 1))+signed(MULTS_1_30(33)(PERCISION) & MULTS_1_30(33)(PERCISION downto 1));
			MULTS_2_15(34)<=signed(MULTS_1_29(34)(PERCISION) & MULTS_1_29(34)(PERCISION downto 1))+signed(MULTS_1_30(34)(PERCISION) & MULTS_1_30(34)(PERCISION downto 1));
			MULTS_2_15(35)<=signed(MULTS_1_29(35)(PERCISION) & MULTS_1_29(35)(PERCISION downto 1))+signed(MULTS_1_30(35)(PERCISION) & MULTS_1_30(35)(PERCISION downto 1));
			MULTS_2_15(36)<=signed(MULTS_1_29(36)(PERCISION) & MULTS_1_29(36)(PERCISION downto 1))+signed(MULTS_1_30(36)(PERCISION) & MULTS_1_30(36)(PERCISION downto 1));
			MULTS_2_15(37)<=signed(MULTS_1_29(37)(PERCISION) & MULTS_1_29(37)(PERCISION downto 1))+signed(MULTS_1_30(37)(PERCISION) & MULTS_1_30(37)(PERCISION downto 1));
			MULTS_2_15(38)<=signed(MULTS_1_29(38)(PERCISION) & MULTS_1_29(38)(PERCISION downto 1))+signed(MULTS_1_30(38)(PERCISION) & MULTS_1_30(38)(PERCISION downto 1));
			MULTS_2_15(39)<=signed(MULTS_1_29(39)(PERCISION) & MULTS_1_29(39)(PERCISION downto 1))+signed(MULTS_1_30(39)(PERCISION) & MULTS_1_30(39)(PERCISION downto 1));
			MULTS_2_15(40)<=signed(MULTS_1_29(40)(PERCISION) & MULTS_1_29(40)(PERCISION downto 1))+signed(MULTS_1_30(40)(PERCISION) & MULTS_1_30(40)(PERCISION downto 1));
			MULTS_2_15(41)<=signed(MULTS_1_29(41)(PERCISION) & MULTS_1_29(41)(PERCISION downto 1))+signed(MULTS_1_30(41)(PERCISION) & MULTS_1_30(41)(PERCISION downto 1));
			MULTS_2_15(42)<=signed(MULTS_1_29(42)(PERCISION) & MULTS_1_29(42)(PERCISION downto 1))+signed(MULTS_1_30(42)(PERCISION) & MULTS_1_30(42)(PERCISION downto 1));
			MULTS_2_15(43)<=signed(MULTS_1_29(43)(PERCISION) & MULTS_1_29(43)(PERCISION downto 1))+signed(MULTS_1_30(43)(PERCISION) & MULTS_1_30(43)(PERCISION downto 1));
			MULTS_2_15(44)<=signed(MULTS_1_29(44)(PERCISION) & MULTS_1_29(44)(PERCISION downto 1))+signed(MULTS_1_30(44)(PERCISION) & MULTS_1_30(44)(PERCISION downto 1));
			MULTS_2_15(45)<=signed(MULTS_1_29(45)(PERCISION) & MULTS_1_29(45)(PERCISION downto 1))+signed(MULTS_1_30(45)(PERCISION) & MULTS_1_30(45)(PERCISION downto 1));
			MULTS_2_15(46)<=signed(MULTS_1_29(46)(PERCISION) & MULTS_1_29(46)(PERCISION downto 1))+signed(MULTS_1_30(46)(PERCISION) & MULTS_1_30(46)(PERCISION downto 1));
			MULTS_2_15(47)<=signed(MULTS_1_29(47)(PERCISION) & MULTS_1_29(47)(PERCISION downto 1))+signed(MULTS_1_30(47)(PERCISION) & MULTS_1_30(47)(PERCISION downto 1));
			MULTS_2_15(48)<=signed(MULTS_1_29(48)(PERCISION) & MULTS_1_29(48)(PERCISION downto 1))+signed(MULTS_1_30(48)(PERCISION) & MULTS_1_30(48)(PERCISION downto 1));
			MULTS_2_15(49)<=signed(MULTS_1_29(49)(PERCISION) & MULTS_1_29(49)(PERCISION downto 1))+signed(MULTS_1_30(49)(PERCISION) & MULTS_1_30(49)(PERCISION downto 1));
			MULTS_2_15(50)<=signed(MULTS_1_29(50)(PERCISION) & MULTS_1_29(50)(PERCISION downto 1))+signed(MULTS_1_30(50)(PERCISION) & MULTS_1_30(50)(PERCISION downto 1));
			MULTS_2_15(51)<=signed(MULTS_1_29(51)(PERCISION) & MULTS_1_29(51)(PERCISION downto 1))+signed(MULTS_1_30(51)(PERCISION) & MULTS_1_30(51)(PERCISION downto 1));
			MULTS_2_15(52)<=signed(MULTS_1_29(52)(PERCISION) & MULTS_1_29(52)(PERCISION downto 1))+signed(MULTS_1_30(52)(PERCISION) & MULTS_1_30(52)(PERCISION downto 1));
			MULTS_2_15(53)<=signed(MULTS_1_29(53)(PERCISION) & MULTS_1_29(53)(PERCISION downto 1))+signed(MULTS_1_30(53)(PERCISION) & MULTS_1_30(53)(PERCISION downto 1));
			MULTS_2_15(54)<=signed(MULTS_1_29(54)(PERCISION) & MULTS_1_29(54)(PERCISION downto 1))+signed(MULTS_1_30(54)(PERCISION) & MULTS_1_30(54)(PERCISION downto 1));
			MULTS_2_15(55)<=signed(MULTS_1_29(55)(PERCISION) & MULTS_1_29(55)(PERCISION downto 1))+signed(MULTS_1_30(55)(PERCISION) & MULTS_1_30(55)(PERCISION downto 1));
			MULTS_2_15(56)<=signed(MULTS_1_29(56)(PERCISION) & MULTS_1_29(56)(PERCISION downto 1))+signed(MULTS_1_30(56)(PERCISION) & MULTS_1_30(56)(PERCISION downto 1));
			MULTS_2_15(57)<=signed(MULTS_1_29(57)(PERCISION) & MULTS_1_29(57)(PERCISION downto 1))+signed(MULTS_1_30(57)(PERCISION) & MULTS_1_30(57)(PERCISION downto 1));
			MULTS_2_15(58)<=signed(MULTS_1_29(58)(PERCISION) & MULTS_1_29(58)(PERCISION downto 1))+signed(MULTS_1_30(58)(PERCISION) & MULTS_1_30(58)(PERCISION downto 1));
			MULTS_2_15(59)<=signed(MULTS_1_29(59)(PERCISION) & MULTS_1_29(59)(PERCISION downto 1))+signed(MULTS_1_30(59)(PERCISION) & MULTS_1_30(59)(PERCISION downto 1));
			MULTS_2_15(60)<=signed(MULTS_1_29(60)(PERCISION) & MULTS_1_29(60)(PERCISION downto 1))+signed(MULTS_1_30(60)(PERCISION) & MULTS_1_30(60)(PERCISION downto 1));
			MULTS_2_15(61)<=signed(MULTS_1_29(61)(PERCISION) & MULTS_1_29(61)(PERCISION downto 1))+signed(MULTS_1_30(61)(PERCISION) & MULTS_1_30(61)(PERCISION downto 1));
			MULTS_2_15(62)<=signed(MULTS_1_29(62)(PERCISION) & MULTS_1_29(62)(PERCISION downto 1))+signed(MULTS_1_30(62)(PERCISION) & MULTS_1_30(62)(PERCISION downto 1));
			MULTS_2_15(63)<=signed(MULTS_1_29(63)(PERCISION) & MULTS_1_29(63)(PERCISION downto 1))+signed(MULTS_1_30(63)(PERCISION) & MULTS_1_30(63)(PERCISION downto 1));
			MULTS_2_15(64)<=signed(MULTS_1_29(64)(PERCISION) & MULTS_1_29(64)(PERCISION downto 1))+signed(MULTS_1_30(64)(PERCISION) & MULTS_1_30(64)(PERCISION downto 1));
			MULTS_2_15(65)<=signed(MULTS_1_29(65)(PERCISION) & MULTS_1_29(65)(PERCISION downto 1))+signed(MULTS_1_30(65)(PERCISION) & MULTS_1_30(65)(PERCISION downto 1));
			MULTS_2_15(66)<=signed(MULTS_1_29(66)(PERCISION) & MULTS_1_29(66)(PERCISION downto 1))+signed(MULTS_1_30(66)(PERCISION) & MULTS_1_30(66)(PERCISION downto 1));
			MULTS_2_15(67)<=signed(MULTS_1_29(67)(PERCISION) & MULTS_1_29(67)(PERCISION downto 1))+signed(MULTS_1_30(67)(PERCISION) & MULTS_1_30(67)(PERCISION downto 1));
			MULTS_2_15(68)<=signed(MULTS_1_29(68)(PERCISION) & MULTS_1_29(68)(PERCISION downto 1))+signed(MULTS_1_30(68)(PERCISION) & MULTS_1_30(68)(PERCISION downto 1));
			MULTS_2_15(69)<=signed(MULTS_1_29(69)(PERCISION) & MULTS_1_29(69)(PERCISION downto 1))+signed(MULTS_1_30(69)(PERCISION) & MULTS_1_30(69)(PERCISION downto 1));
			MULTS_2_15(70)<=signed(MULTS_1_29(70)(PERCISION) & MULTS_1_29(70)(PERCISION downto 1))+signed(MULTS_1_30(70)(PERCISION) & MULTS_1_30(70)(PERCISION downto 1));
			MULTS_2_15(71)<=signed(MULTS_1_29(71)(PERCISION) & MULTS_1_29(71)(PERCISION downto 1))+signed(MULTS_1_30(71)(PERCISION) & MULTS_1_30(71)(PERCISION downto 1));
			MULTS_2_15(72)<=signed(MULTS_1_29(72)(PERCISION) & MULTS_1_29(72)(PERCISION downto 1))+signed(MULTS_1_30(72)(PERCISION) & MULTS_1_30(72)(PERCISION downto 1));
			MULTS_2_15(73)<=signed(MULTS_1_29(73)(PERCISION) & MULTS_1_29(73)(PERCISION downto 1))+signed(MULTS_1_30(73)(PERCISION) & MULTS_1_30(73)(PERCISION downto 1));
			MULTS_2_15(74)<=signed(MULTS_1_29(74)(PERCISION) & MULTS_1_29(74)(PERCISION downto 1))+signed(MULTS_1_30(74)(PERCISION) & MULTS_1_30(74)(PERCISION downto 1));
			MULTS_2_15(75)<=signed(MULTS_1_29(75)(PERCISION) & MULTS_1_29(75)(PERCISION downto 1))+signed(MULTS_1_30(75)(PERCISION) & MULTS_1_30(75)(PERCISION downto 1));
			MULTS_2_15(76)<=signed(MULTS_1_29(76)(PERCISION) & MULTS_1_29(76)(PERCISION downto 1))+signed(MULTS_1_30(76)(PERCISION) & MULTS_1_30(76)(PERCISION downto 1));
			MULTS_2_15(77)<=signed(MULTS_1_29(77)(PERCISION) & MULTS_1_29(77)(PERCISION downto 1))+signed(MULTS_1_30(77)(PERCISION) & MULTS_1_30(77)(PERCISION downto 1));
			MULTS_2_15(78)<=signed(MULTS_1_29(78)(PERCISION) & MULTS_1_29(78)(PERCISION downto 1))+signed(MULTS_1_30(78)(PERCISION) & MULTS_1_30(78)(PERCISION downto 1));
			MULTS_2_15(79)<=signed(MULTS_1_29(79)(PERCISION) & MULTS_1_29(79)(PERCISION downto 1))+signed(MULTS_1_30(79)(PERCISION) & MULTS_1_30(79)(PERCISION downto 1));
			MULTS_2_15(80)<=signed(MULTS_1_29(80)(PERCISION) & MULTS_1_29(80)(PERCISION downto 1))+signed(MULTS_1_30(80)(PERCISION) & MULTS_1_30(80)(PERCISION downto 1));
			MULTS_2_15(81)<=signed(MULTS_1_29(81)(PERCISION) & MULTS_1_29(81)(PERCISION downto 1))+signed(MULTS_1_30(81)(PERCISION) & MULTS_1_30(81)(PERCISION downto 1));
			MULTS_2_15(82)<=signed(MULTS_1_29(82)(PERCISION) & MULTS_1_29(82)(PERCISION downto 1))+signed(MULTS_1_30(82)(PERCISION) & MULTS_1_30(82)(PERCISION downto 1));
			MULTS_2_15(83)<=signed(MULTS_1_29(83)(PERCISION) & MULTS_1_29(83)(PERCISION downto 1))+signed(MULTS_1_30(83)(PERCISION) & MULTS_1_30(83)(PERCISION downto 1));



                         EN_SUM_MULT_3<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_3 = '1' then
			------------------------------------STAGE-3--------------------------------------
			MULTS_3_1(0)<=signed(MULTS_2_1(0)(PERCISION) & MULTS_2_1(0)(PERCISION downto 1))+signed(MULTS_2_2(0)(PERCISION) & MULTS_2_2(0)(PERCISION downto 1));
			MULTS_3_1(1)<=signed(MULTS_2_1(1)(PERCISION) & MULTS_2_1(1)(PERCISION downto 1))+signed(MULTS_2_2(1)(PERCISION) & MULTS_2_2(1)(PERCISION downto 1));
			MULTS_3_1(2)<=signed(MULTS_2_1(2)(PERCISION) & MULTS_2_1(2)(PERCISION downto 1))+signed(MULTS_2_2(2)(PERCISION) & MULTS_2_2(2)(PERCISION downto 1));
			MULTS_3_1(3)<=signed(MULTS_2_1(3)(PERCISION) & MULTS_2_1(3)(PERCISION downto 1))+signed(MULTS_2_2(3)(PERCISION) & MULTS_2_2(3)(PERCISION downto 1));
			MULTS_3_1(4)<=signed(MULTS_2_1(4)(PERCISION) & MULTS_2_1(4)(PERCISION downto 1))+signed(MULTS_2_2(4)(PERCISION) & MULTS_2_2(4)(PERCISION downto 1));
			MULTS_3_1(5)<=signed(MULTS_2_1(5)(PERCISION) & MULTS_2_1(5)(PERCISION downto 1))+signed(MULTS_2_2(5)(PERCISION) & MULTS_2_2(5)(PERCISION downto 1));
			MULTS_3_1(6)<=signed(MULTS_2_1(6)(PERCISION) & MULTS_2_1(6)(PERCISION downto 1))+signed(MULTS_2_2(6)(PERCISION) & MULTS_2_2(6)(PERCISION downto 1));
			MULTS_3_1(7)<=signed(MULTS_2_1(7)(PERCISION) & MULTS_2_1(7)(PERCISION downto 1))+signed(MULTS_2_2(7)(PERCISION) & MULTS_2_2(7)(PERCISION downto 1));
			MULTS_3_1(8)<=signed(MULTS_2_1(8)(PERCISION) & MULTS_2_1(8)(PERCISION downto 1))+signed(MULTS_2_2(8)(PERCISION) & MULTS_2_2(8)(PERCISION downto 1));
			MULTS_3_1(9)<=signed(MULTS_2_1(9)(PERCISION) & MULTS_2_1(9)(PERCISION downto 1))+signed(MULTS_2_2(9)(PERCISION) & MULTS_2_2(9)(PERCISION downto 1));
			MULTS_3_1(10)<=signed(MULTS_2_1(10)(PERCISION) & MULTS_2_1(10)(PERCISION downto 1))+signed(MULTS_2_2(10)(PERCISION) & MULTS_2_2(10)(PERCISION downto 1));
			MULTS_3_1(11)<=signed(MULTS_2_1(11)(PERCISION) & MULTS_2_1(11)(PERCISION downto 1))+signed(MULTS_2_2(11)(PERCISION) & MULTS_2_2(11)(PERCISION downto 1));
			MULTS_3_1(12)<=signed(MULTS_2_1(12)(PERCISION) & MULTS_2_1(12)(PERCISION downto 1))+signed(MULTS_2_2(12)(PERCISION) & MULTS_2_2(12)(PERCISION downto 1));
			MULTS_3_1(13)<=signed(MULTS_2_1(13)(PERCISION) & MULTS_2_1(13)(PERCISION downto 1))+signed(MULTS_2_2(13)(PERCISION) & MULTS_2_2(13)(PERCISION downto 1));
			MULTS_3_1(14)<=signed(MULTS_2_1(14)(PERCISION) & MULTS_2_1(14)(PERCISION downto 1))+signed(MULTS_2_2(14)(PERCISION) & MULTS_2_2(14)(PERCISION downto 1));
			MULTS_3_1(15)<=signed(MULTS_2_1(15)(PERCISION) & MULTS_2_1(15)(PERCISION downto 1))+signed(MULTS_2_2(15)(PERCISION) & MULTS_2_2(15)(PERCISION downto 1));
			MULTS_3_1(16)<=signed(MULTS_2_1(16)(PERCISION) & MULTS_2_1(16)(PERCISION downto 1))+signed(MULTS_2_2(16)(PERCISION) & MULTS_2_2(16)(PERCISION downto 1));
			MULTS_3_1(17)<=signed(MULTS_2_1(17)(PERCISION) & MULTS_2_1(17)(PERCISION downto 1))+signed(MULTS_2_2(17)(PERCISION) & MULTS_2_2(17)(PERCISION downto 1));
			MULTS_3_1(18)<=signed(MULTS_2_1(18)(PERCISION) & MULTS_2_1(18)(PERCISION downto 1))+signed(MULTS_2_2(18)(PERCISION) & MULTS_2_2(18)(PERCISION downto 1));
			MULTS_3_1(19)<=signed(MULTS_2_1(19)(PERCISION) & MULTS_2_1(19)(PERCISION downto 1))+signed(MULTS_2_2(19)(PERCISION) & MULTS_2_2(19)(PERCISION downto 1));
			MULTS_3_1(20)<=signed(MULTS_2_1(20)(PERCISION) & MULTS_2_1(20)(PERCISION downto 1))+signed(MULTS_2_2(20)(PERCISION) & MULTS_2_2(20)(PERCISION downto 1));
			MULTS_3_1(21)<=signed(MULTS_2_1(21)(PERCISION) & MULTS_2_1(21)(PERCISION downto 1))+signed(MULTS_2_2(21)(PERCISION) & MULTS_2_2(21)(PERCISION downto 1));
			MULTS_3_1(22)<=signed(MULTS_2_1(22)(PERCISION) & MULTS_2_1(22)(PERCISION downto 1))+signed(MULTS_2_2(22)(PERCISION) & MULTS_2_2(22)(PERCISION downto 1));
			MULTS_3_1(23)<=signed(MULTS_2_1(23)(PERCISION) & MULTS_2_1(23)(PERCISION downto 1))+signed(MULTS_2_2(23)(PERCISION) & MULTS_2_2(23)(PERCISION downto 1));
			MULTS_3_1(24)<=signed(MULTS_2_1(24)(PERCISION) & MULTS_2_1(24)(PERCISION downto 1))+signed(MULTS_2_2(24)(PERCISION) & MULTS_2_2(24)(PERCISION downto 1));
			MULTS_3_1(25)<=signed(MULTS_2_1(25)(PERCISION) & MULTS_2_1(25)(PERCISION downto 1))+signed(MULTS_2_2(25)(PERCISION) & MULTS_2_2(25)(PERCISION downto 1));
			MULTS_3_1(26)<=signed(MULTS_2_1(26)(PERCISION) & MULTS_2_1(26)(PERCISION downto 1))+signed(MULTS_2_2(26)(PERCISION) & MULTS_2_2(26)(PERCISION downto 1));
			MULTS_3_1(27)<=signed(MULTS_2_1(27)(PERCISION) & MULTS_2_1(27)(PERCISION downto 1))+signed(MULTS_2_2(27)(PERCISION) & MULTS_2_2(27)(PERCISION downto 1));
			MULTS_3_1(28)<=signed(MULTS_2_1(28)(PERCISION) & MULTS_2_1(28)(PERCISION downto 1))+signed(MULTS_2_2(28)(PERCISION) & MULTS_2_2(28)(PERCISION downto 1));
			MULTS_3_1(29)<=signed(MULTS_2_1(29)(PERCISION) & MULTS_2_1(29)(PERCISION downto 1))+signed(MULTS_2_2(29)(PERCISION) & MULTS_2_2(29)(PERCISION downto 1));
			MULTS_3_1(30)<=signed(MULTS_2_1(30)(PERCISION) & MULTS_2_1(30)(PERCISION downto 1))+signed(MULTS_2_2(30)(PERCISION) & MULTS_2_2(30)(PERCISION downto 1));
			MULTS_3_1(31)<=signed(MULTS_2_1(31)(PERCISION) & MULTS_2_1(31)(PERCISION downto 1))+signed(MULTS_2_2(31)(PERCISION) & MULTS_2_2(31)(PERCISION downto 1));
			MULTS_3_1(32)<=signed(MULTS_2_1(32)(PERCISION) & MULTS_2_1(32)(PERCISION downto 1))+signed(MULTS_2_2(32)(PERCISION) & MULTS_2_2(32)(PERCISION downto 1));
			MULTS_3_1(33)<=signed(MULTS_2_1(33)(PERCISION) & MULTS_2_1(33)(PERCISION downto 1))+signed(MULTS_2_2(33)(PERCISION) & MULTS_2_2(33)(PERCISION downto 1));
			MULTS_3_1(34)<=signed(MULTS_2_1(34)(PERCISION) & MULTS_2_1(34)(PERCISION downto 1))+signed(MULTS_2_2(34)(PERCISION) & MULTS_2_2(34)(PERCISION downto 1));
			MULTS_3_1(35)<=signed(MULTS_2_1(35)(PERCISION) & MULTS_2_1(35)(PERCISION downto 1))+signed(MULTS_2_2(35)(PERCISION) & MULTS_2_2(35)(PERCISION downto 1));
			MULTS_3_1(36)<=signed(MULTS_2_1(36)(PERCISION) & MULTS_2_1(36)(PERCISION downto 1))+signed(MULTS_2_2(36)(PERCISION) & MULTS_2_2(36)(PERCISION downto 1));
			MULTS_3_1(37)<=signed(MULTS_2_1(37)(PERCISION) & MULTS_2_1(37)(PERCISION downto 1))+signed(MULTS_2_2(37)(PERCISION) & MULTS_2_2(37)(PERCISION downto 1));
			MULTS_3_1(38)<=signed(MULTS_2_1(38)(PERCISION) & MULTS_2_1(38)(PERCISION downto 1))+signed(MULTS_2_2(38)(PERCISION) & MULTS_2_2(38)(PERCISION downto 1));
			MULTS_3_1(39)<=signed(MULTS_2_1(39)(PERCISION) & MULTS_2_1(39)(PERCISION downto 1))+signed(MULTS_2_2(39)(PERCISION) & MULTS_2_2(39)(PERCISION downto 1));
			MULTS_3_1(40)<=signed(MULTS_2_1(40)(PERCISION) & MULTS_2_1(40)(PERCISION downto 1))+signed(MULTS_2_2(40)(PERCISION) & MULTS_2_2(40)(PERCISION downto 1));
			MULTS_3_1(41)<=signed(MULTS_2_1(41)(PERCISION) & MULTS_2_1(41)(PERCISION downto 1))+signed(MULTS_2_2(41)(PERCISION) & MULTS_2_2(41)(PERCISION downto 1));
			MULTS_3_1(42)<=signed(MULTS_2_1(42)(PERCISION) & MULTS_2_1(42)(PERCISION downto 1))+signed(MULTS_2_2(42)(PERCISION) & MULTS_2_2(42)(PERCISION downto 1));
			MULTS_3_1(43)<=signed(MULTS_2_1(43)(PERCISION) & MULTS_2_1(43)(PERCISION downto 1))+signed(MULTS_2_2(43)(PERCISION) & MULTS_2_2(43)(PERCISION downto 1));
			MULTS_3_1(44)<=signed(MULTS_2_1(44)(PERCISION) & MULTS_2_1(44)(PERCISION downto 1))+signed(MULTS_2_2(44)(PERCISION) & MULTS_2_2(44)(PERCISION downto 1));
			MULTS_3_1(45)<=signed(MULTS_2_1(45)(PERCISION) & MULTS_2_1(45)(PERCISION downto 1))+signed(MULTS_2_2(45)(PERCISION) & MULTS_2_2(45)(PERCISION downto 1));
			MULTS_3_1(46)<=signed(MULTS_2_1(46)(PERCISION) & MULTS_2_1(46)(PERCISION downto 1))+signed(MULTS_2_2(46)(PERCISION) & MULTS_2_2(46)(PERCISION downto 1));
			MULTS_3_1(47)<=signed(MULTS_2_1(47)(PERCISION) & MULTS_2_1(47)(PERCISION downto 1))+signed(MULTS_2_2(47)(PERCISION) & MULTS_2_2(47)(PERCISION downto 1));
			MULTS_3_1(48)<=signed(MULTS_2_1(48)(PERCISION) & MULTS_2_1(48)(PERCISION downto 1))+signed(MULTS_2_2(48)(PERCISION) & MULTS_2_2(48)(PERCISION downto 1));
			MULTS_3_1(49)<=signed(MULTS_2_1(49)(PERCISION) & MULTS_2_1(49)(PERCISION downto 1))+signed(MULTS_2_2(49)(PERCISION) & MULTS_2_2(49)(PERCISION downto 1));
			MULTS_3_1(50)<=signed(MULTS_2_1(50)(PERCISION) & MULTS_2_1(50)(PERCISION downto 1))+signed(MULTS_2_2(50)(PERCISION) & MULTS_2_2(50)(PERCISION downto 1));
			MULTS_3_1(51)<=signed(MULTS_2_1(51)(PERCISION) & MULTS_2_1(51)(PERCISION downto 1))+signed(MULTS_2_2(51)(PERCISION) & MULTS_2_2(51)(PERCISION downto 1));
			MULTS_3_1(52)<=signed(MULTS_2_1(52)(PERCISION) & MULTS_2_1(52)(PERCISION downto 1))+signed(MULTS_2_2(52)(PERCISION) & MULTS_2_2(52)(PERCISION downto 1));
			MULTS_3_1(53)<=signed(MULTS_2_1(53)(PERCISION) & MULTS_2_1(53)(PERCISION downto 1))+signed(MULTS_2_2(53)(PERCISION) & MULTS_2_2(53)(PERCISION downto 1));
			MULTS_3_1(54)<=signed(MULTS_2_1(54)(PERCISION) & MULTS_2_1(54)(PERCISION downto 1))+signed(MULTS_2_2(54)(PERCISION) & MULTS_2_2(54)(PERCISION downto 1));
			MULTS_3_1(55)<=signed(MULTS_2_1(55)(PERCISION) & MULTS_2_1(55)(PERCISION downto 1))+signed(MULTS_2_2(55)(PERCISION) & MULTS_2_2(55)(PERCISION downto 1));
			MULTS_3_1(56)<=signed(MULTS_2_1(56)(PERCISION) & MULTS_2_1(56)(PERCISION downto 1))+signed(MULTS_2_2(56)(PERCISION) & MULTS_2_2(56)(PERCISION downto 1));
			MULTS_3_1(57)<=signed(MULTS_2_1(57)(PERCISION) & MULTS_2_1(57)(PERCISION downto 1))+signed(MULTS_2_2(57)(PERCISION) & MULTS_2_2(57)(PERCISION downto 1));
			MULTS_3_1(58)<=signed(MULTS_2_1(58)(PERCISION) & MULTS_2_1(58)(PERCISION downto 1))+signed(MULTS_2_2(58)(PERCISION) & MULTS_2_2(58)(PERCISION downto 1));
			MULTS_3_1(59)<=signed(MULTS_2_1(59)(PERCISION) & MULTS_2_1(59)(PERCISION downto 1))+signed(MULTS_2_2(59)(PERCISION) & MULTS_2_2(59)(PERCISION downto 1));
			MULTS_3_1(60)<=signed(MULTS_2_1(60)(PERCISION) & MULTS_2_1(60)(PERCISION downto 1))+signed(MULTS_2_2(60)(PERCISION) & MULTS_2_2(60)(PERCISION downto 1));
			MULTS_3_1(61)<=signed(MULTS_2_1(61)(PERCISION) & MULTS_2_1(61)(PERCISION downto 1))+signed(MULTS_2_2(61)(PERCISION) & MULTS_2_2(61)(PERCISION downto 1));
			MULTS_3_1(62)<=signed(MULTS_2_1(62)(PERCISION) & MULTS_2_1(62)(PERCISION downto 1))+signed(MULTS_2_2(62)(PERCISION) & MULTS_2_2(62)(PERCISION downto 1));
			MULTS_3_1(63)<=signed(MULTS_2_1(63)(PERCISION) & MULTS_2_1(63)(PERCISION downto 1))+signed(MULTS_2_2(63)(PERCISION) & MULTS_2_2(63)(PERCISION downto 1));
			MULTS_3_1(64)<=signed(MULTS_2_1(64)(PERCISION) & MULTS_2_1(64)(PERCISION downto 1))+signed(MULTS_2_2(64)(PERCISION) & MULTS_2_2(64)(PERCISION downto 1));
			MULTS_3_1(65)<=signed(MULTS_2_1(65)(PERCISION) & MULTS_2_1(65)(PERCISION downto 1))+signed(MULTS_2_2(65)(PERCISION) & MULTS_2_2(65)(PERCISION downto 1));
			MULTS_3_1(66)<=signed(MULTS_2_1(66)(PERCISION) & MULTS_2_1(66)(PERCISION downto 1))+signed(MULTS_2_2(66)(PERCISION) & MULTS_2_2(66)(PERCISION downto 1));
			MULTS_3_1(67)<=signed(MULTS_2_1(67)(PERCISION) & MULTS_2_1(67)(PERCISION downto 1))+signed(MULTS_2_2(67)(PERCISION) & MULTS_2_2(67)(PERCISION downto 1));
			MULTS_3_1(68)<=signed(MULTS_2_1(68)(PERCISION) & MULTS_2_1(68)(PERCISION downto 1))+signed(MULTS_2_2(68)(PERCISION) & MULTS_2_2(68)(PERCISION downto 1));
			MULTS_3_1(69)<=signed(MULTS_2_1(69)(PERCISION) & MULTS_2_1(69)(PERCISION downto 1))+signed(MULTS_2_2(69)(PERCISION) & MULTS_2_2(69)(PERCISION downto 1));
			MULTS_3_1(70)<=signed(MULTS_2_1(70)(PERCISION) & MULTS_2_1(70)(PERCISION downto 1))+signed(MULTS_2_2(70)(PERCISION) & MULTS_2_2(70)(PERCISION downto 1));
			MULTS_3_1(71)<=signed(MULTS_2_1(71)(PERCISION) & MULTS_2_1(71)(PERCISION downto 1))+signed(MULTS_2_2(71)(PERCISION) & MULTS_2_2(71)(PERCISION downto 1));
			MULTS_3_1(72)<=signed(MULTS_2_1(72)(PERCISION) & MULTS_2_1(72)(PERCISION downto 1))+signed(MULTS_2_2(72)(PERCISION) & MULTS_2_2(72)(PERCISION downto 1));
			MULTS_3_1(73)<=signed(MULTS_2_1(73)(PERCISION) & MULTS_2_1(73)(PERCISION downto 1))+signed(MULTS_2_2(73)(PERCISION) & MULTS_2_2(73)(PERCISION downto 1));
			MULTS_3_1(74)<=signed(MULTS_2_1(74)(PERCISION) & MULTS_2_1(74)(PERCISION downto 1))+signed(MULTS_2_2(74)(PERCISION) & MULTS_2_2(74)(PERCISION downto 1));
			MULTS_3_1(75)<=signed(MULTS_2_1(75)(PERCISION) & MULTS_2_1(75)(PERCISION downto 1))+signed(MULTS_2_2(75)(PERCISION) & MULTS_2_2(75)(PERCISION downto 1));
			MULTS_3_1(76)<=signed(MULTS_2_1(76)(PERCISION) & MULTS_2_1(76)(PERCISION downto 1))+signed(MULTS_2_2(76)(PERCISION) & MULTS_2_2(76)(PERCISION downto 1));
			MULTS_3_1(77)<=signed(MULTS_2_1(77)(PERCISION) & MULTS_2_1(77)(PERCISION downto 1))+signed(MULTS_2_2(77)(PERCISION) & MULTS_2_2(77)(PERCISION downto 1));
			MULTS_3_1(78)<=signed(MULTS_2_1(78)(PERCISION) & MULTS_2_1(78)(PERCISION downto 1))+signed(MULTS_2_2(78)(PERCISION) & MULTS_2_2(78)(PERCISION downto 1));
			MULTS_3_1(79)<=signed(MULTS_2_1(79)(PERCISION) & MULTS_2_1(79)(PERCISION downto 1))+signed(MULTS_2_2(79)(PERCISION) & MULTS_2_2(79)(PERCISION downto 1));
			MULTS_3_1(80)<=signed(MULTS_2_1(80)(PERCISION) & MULTS_2_1(80)(PERCISION downto 1))+signed(MULTS_2_2(80)(PERCISION) & MULTS_2_2(80)(PERCISION downto 1));
			MULTS_3_1(81)<=signed(MULTS_2_1(81)(PERCISION) & MULTS_2_1(81)(PERCISION downto 1))+signed(MULTS_2_2(81)(PERCISION) & MULTS_2_2(81)(PERCISION downto 1));
			MULTS_3_1(82)<=signed(MULTS_2_1(82)(PERCISION) & MULTS_2_1(82)(PERCISION downto 1))+signed(MULTS_2_2(82)(PERCISION) & MULTS_2_2(82)(PERCISION downto 1));
			MULTS_3_1(83)<=signed(MULTS_2_1(83)(PERCISION) & MULTS_2_1(83)(PERCISION downto 1))+signed(MULTS_2_2(83)(PERCISION) & MULTS_2_2(83)(PERCISION downto 1));

			MULTS_3_2(0)<=signed(MULTS_2_3(0)(PERCISION) & MULTS_2_3(0)(PERCISION downto 1))+signed(MULTS_2_4(0)(PERCISION) & MULTS_2_4(0)(PERCISION downto 1));
			MULTS_3_2(1)<=signed(MULTS_2_3(1)(PERCISION) & MULTS_2_3(1)(PERCISION downto 1))+signed(MULTS_2_4(1)(PERCISION) & MULTS_2_4(1)(PERCISION downto 1));
			MULTS_3_2(2)<=signed(MULTS_2_3(2)(PERCISION) & MULTS_2_3(2)(PERCISION downto 1))+signed(MULTS_2_4(2)(PERCISION) & MULTS_2_4(2)(PERCISION downto 1));
			MULTS_3_2(3)<=signed(MULTS_2_3(3)(PERCISION) & MULTS_2_3(3)(PERCISION downto 1))+signed(MULTS_2_4(3)(PERCISION) & MULTS_2_4(3)(PERCISION downto 1));
			MULTS_3_2(4)<=signed(MULTS_2_3(4)(PERCISION) & MULTS_2_3(4)(PERCISION downto 1))+signed(MULTS_2_4(4)(PERCISION) & MULTS_2_4(4)(PERCISION downto 1));
			MULTS_3_2(5)<=signed(MULTS_2_3(5)(PERCISION) & MULTS_2_3(5)(PERCISION downto 1))+signed(MULTS_2_4(5)(PERCISION) & MULTS_2_4(5)(PERCISION downto 1));
			MULTS_3_2(6)<=signed(MULTS_2_3(6)(PERCISION) & MULTS_2_3(6)(PERCISION downto 1))+signed(MULTS_2_4(6)(PERCISION) & MULTS_2_4(6)(PERCISION downto 1));
			MULTS_3_2(7)<=signed(MULTS_2_3(7)(PERCISION) & MULTS_2_3(7)(PERCISION downto 1))+signed(MULTS_2_4(7)(PERCISION) & MULTS_2_4(7)(PERCISION downto 1));
			MULTS_3_2(8)<=signed(MULTS_2_3(8)(PERCISION) & MULTS_2_3(8)(PERCISION downto 1))+signed(MULTS_2_4(8)(PERCISION) & MULTS_2_4(8)(PERCISION downto 1));
			MULTS_3_2(9)<=signed(MULTS_2_3(9)(PERCISION) & MULTS_2_3(9)(PERCISION downto 1))+signed(MULTS_2_4(9)(PERCISION) & MULTS_2_4(9)(PERCISION downto 1));
			MULTS_3_2(10)<=signed(MULTS_2_3(10)(PERCISION) & MULTS_2_3(10)(PERCISION downto 1))+signed(MULTS_2_4(10)(PERCISION) & MULTS_2_4(10)(PERCISION downto 1));
			MULTS_3_2(11)<=signed(MULTS_2_3(11)(PERCISION) & MULTS_2_3(11)(PERCISION downto 1))+signed(MULTS_2_4(11)(PERCISION) & MULTS_2_4(11)(PERCISION downto 1));
			MULTS_3_2(12)<=signed(MULTS_2_3(12)(PERCISION) & MULTS_2_3(12)(PERCISION downto 1))+signed(MULTS_2_4(12)(PERCISION) & MULTS_2_4(12)(PERCISION downto 1));
			MULTS_3_2(13)<=signed(MULTS_2_3(13)(PERCISION) & MULTS_2_3(13)(PERCISION downto 1))+signed(MULTS_2_4(13)(PERCISION) & MULTS_2_4(13)(PERCISION downto 1));
			MULTS_3_2(14)<=signed(MULTS_2_3(14)(PERCISION) & MULTS_2_3(14)(PERCISION downto 1))+signed(MULTS_2_4(14)(PERCISION) & MULTS_2_4(14)(PERCISION downto 1));
			MULTS_3_2(15)<=signed(MULTS_2_3(15)(PERCISION) & MULTS_2_3(15)(PERCISION downto 1))+signed(MULTS_2_4(15)(PERCISION) & MULTS_2_4(15)(PERCISION downto 1));
			MULTS_3_2(16)<=signed(MULTS_2_3(16)(PERCISION) & MULTS_2_3(16)(PERCISION downto 1))+signed(MULTS_2_4(16)(PERCISION) & MULTS_2_4(16)(PERCISION downto 1));
			MULTS_3_2(17)<=signed(MULTS_2_3(17)(PERCISION) & MULTS_2_3(17)(PERCISION downto 1))+signed(MULTS_2_4(17)(PERCISION) & MULTS_2_4(17)(PERCISION downto 1));
			MULTS_3_2(18)<=signed(MULTS_2_3(18)(PERCISION) & MULTS_2_3(18)(PERCISION downto 1))+signed(MULTS_2_4(18)(PERCISION) & MULTS_2_4(18)(PERCISION downto 1));
			MULTS_3_2(19)<=signed(MULTS_2_3(19)(PERCISION) & MULTS_2_3(19)(PERCISION downto 1))+signed(MULTS_2_4(19)(PERCISION) & MULTS_2_4(19)(PERCISION downto 1));
			MULTS_3_2(20)<=signed(MULTS_2_3(20)(PERCISION) & MULTS_2_3(20)(PERCISION downto 1))+signed(MULTS_2_4(20)(PERCISION) & MULTS_2_4(20)(PERCISION downto 1));
			MULTS_3_2(21)<=signed(MULTS_2_3(21)(PERCISION) & MULTS_2_3(21)(PERCISION downto 1))+signed(MULTS_2_4(21)(PERCISION) & MULTS_2_4(21)(PERCISION downto 1));
			MULTS_3_2(22)<=signed(MULTS_2_3(22)(PERCISION) & MULTS_2_3(22)(PERCISION downto 1))+signed(MULTS_2_4(22)(PERCISION) & MULTS_2_4(22)(PERCISION downto 1));
			MULTS_3_2(23)<=signed(MULTS_2_3(23)(PERCISION) & MULTS_2_3(23)(PERCISION downto 1))+signed(MULTS_2_4(23)(PERCISION) & MULTS_2_4(23)(PERCISION downto 1));
			MULTS_3_2(24)<=signed(MULTS_2_3(24)(PERCISION) & MULTS_2_3(24)(PERCISION downto 1))+signed(MULTS_2_4(24)(PERCISION) & MULTS_2_4(24)(PERCISION downto 1));
			MULTS_3_2(25)<=signed(MULTS_2_3(25)(PERCISION) & MULTS_2_3(25)(PERCISION downto 1))+signed(MULTS_2_4(25)(PERCISION) & MULTS_2_4(25)(PERCISION downto 1));
			MULTS_3_2(26)<=signed(MULTS_2_3(26)(PERCISION) & MULTS_2_3(26)(PERCISION downto 1))+signed(MULTS_2_4(26)(PERCISION) & MULTS_2_4(26)(PERCISION downto 1));
			MULTS_3_2(27)<=signed(MULTS_2_3(27)(PERCISION) & MULTS_2_3(27)(PERCISION downto 1))+signed(MULTS_2_4(27)(PERCISION) & MULTS_2_4(27)(PERCISION downto 1));
			MULTS_3_2(28)<=signed(MULTS_2_3(28)(PERCISION) & MULTS_2_3(28)(PERCISION downto 1))+signed(MULTS_2_4(28)(PERCISION) & MULTS_2_4(28)(PERCISION downto 1));
			MULTS_3_2(29)<=signed(MULTS_2_3(29)(PERCISION) & MULTS_2_3(29)(PERCISION downto 1))+signed(MULTS_2_4(29)(PERCISION) & MULTS_2_4(29)(PERCISION downto 1));
			MULTS_3_2(30)<=signed(MULTS_2_3(30)(PERCISION) & MULTS_2_3(30)(PERCISION downto 1))+signed(MULTS_2_4(30)(PERCISION) & MULTS_2_4(30)(PERCISION downto 1));
			MULTS_3_2(31)<=signed(MULTS_2_3(31)(PERCISION) & MULTS_2_3(31)(PERCISION downto 1))+signed(MULTS_2_4(31)(PERCISION) & MULTS_2_4(31)(PERCISION downto 1));
			MULTS_3_2(32)<=signed(MULTS_2_3(32)(PERCISION) & MULTS_2_3(32)(PERCISION downto 1))+signed(MULTS_2_4(32)(PERCISION) & MULTS_2_4(32)(PERCISION downto 1));
			MULTS_3_2(33)<=signed(MULTS_2_3(33)(PERCISION) & MULTS_2_3(33)(PERCISION downto 1))+signed(MULTS_2_4(33)(PERCISION) & MULTS_2_4(33)(PERCISION downto 1));
			MULTS_3_2(34)<=signed(MULTS_2_3(34)(PERCISION) & MULTS_2_3(34)(PERCISION downto 1))+signed(MULTS_2_4(34)(PERCISION) & MULTS_2_4(34)(PERCISION downto 1));
			MULTS_3_2(35)<=signed(MULTS_2_3(35)(PERCISION) & MULTS_2_3(35)(PERCISION downto 1))+signed(MULTS_2_4(35)(PERCISION) & MULTS_2_4(35)(PERCISION downto 1));
			MULTS_3_2(36)<=signed(MULTS_2_3(36)(PERCISION) & MULTS_2_3(36)(PERCISION downto 1))+signed(MULTS_2_4(36)(PERCISION) & MULTS_2_4(36)(PERCISION downto 1));
			MULTS_3_2(37)<=signed(MULTS_2_3(37)(PERCISION) & MULTS_2_3(37)(PERCISION downto 1))+signed(MULTS_2_4(37)(PERCISION) & MULTS_2_4(37)(PERCISION downto 1));
			MULTS_3_2(38)<=signed(MULTS_2_3(38)(PERCISION) & MULTS_2_3(38)(PERCISION downto 1))+signed(MULTS_2_4(38)(PERCISION) & MULTS_2_4(38)(PERCISION downto 1));
			MULTS_3_2(39)<=signed(MULTS_2_3(39)(PERCISION) & MULTS_2_3(39)(PERCISION downto 1))+signed(MULTS_2_4(39)(PERCISION) & MULTS_2_4(39)(PERCISION downto 1));
			MULTS_3_2(40)<=signed(MULTS_2_3(40)(PERCISION) & MULTS_2_3(40)(PERCISION downto 1))+signed(MULTS_2_4(40)(PERCISION) & MULTS_2_4(40)(PERCISION downto 1));
			MULTS_3_2(41)<=signed(MULTS_2_3(41)(PERCISION) & MULTS_2_3(41)(PERCISION downto 1))+signed(MULTS_2_4(41)(PERCISION) & MULTS_2_4(41)(PERCISION downto 1));
			MULTS_3_2(42)<=signed(MULTS_2_3(42)(PERCISION) & MULTS_2_3(42)(PERCISION downto 1))+signed(MULTS_2_4(42)(PERCISION) & MULTS_2_4(42)(PERCISION downto 1));
			MULTS_3_2(43)<=signed(MULTS_2_3(43)(PERCISION) & MULTS_2_3(43)(PERCISION downto 1))+signed(MULTS_2_4(43)(PERCISION) & MULTS_2_4(43)(PERCISION downto 1));
			MULTS_3_2(44)<=signed(MULTS_2_3(44)(PERCISION) & MULTS_2_3(44)(PERCISION downto 1))+signed(MULTS_2_4(44)(PERCISION) & MULTS_2_4(44)(PERCISION downto 1));
			MULTS_3_2(45)<=signed(MULTS_2_3(45)(PERCISION) & MULTS_2_3(45)(PERCISION downto 1))+signed(MULTS_2_4(45)(PERCISION) & MULTS_2_4(45)(PERCISION downto 1));
			MULTS_3_2(46)<=signed(MULTS_2_3(46)(PERCISION) & MULTS_2_3(46)(PERCISION downto 1))+signed(MULTS_2_4(46)(PERCISION) & MULTS_2_4(46)(PERCISION downto 1));
			MULTS_3_2(47)<=signed(MULTS_2_3(47)(PERCISION) & MULTS_2_3(47)(PERCISION downto 1))+signed(MULTS_2_4(47)(PERCISION) & MULTS_2_4(47)(PERCISION downto 1));
			MULTS_3_2(48)<=signed(MULTS_2_3(48)(PERCISION) & MULTS_2_3(48)(PERCISION downto 1))+signed(MULTS_2_4(48)(PERCISION) & MULTS_2_4(48)(PERCISION downto 1));
			MULTS_3_2(49)<=signed(MULTS_2_3(49)(PERCISION) & MULTS_2_3(49)(PERCISION downto 1))+signed(MULTS_2_4(49)(PERCISION) & MULTS_2_4(49)(PERCISION downto 1));
			MULTS_3_2(50)<=signed(MULTS_2_3(50)(PERCISION) & MULTS_2_3(50)(PERCISION downto 1))+signed(MULTS_2_4(50)(PERCISION) & MULTS_2_4(50)(PERCISION downto 1));
			MULTS_3_2(51)<=signed(MULTS_2_3(51)(PERCISION) & MULTS_2_3(51)(PERCISION downto 1))+signed(MULTS_2_4(51)(PERCISION) & MULTS_2_4(51)(PERCISION downto 1));
			MULTS_3_2(52)<=signed(MULTS_2_3(52)(PERCISION) & MULTS_2_3(52)(PERCISION downto 1))+signed(MULTS_2_4(52)(PERCISION) & MULTS_2_4(52)(PERCISION downto 1));
			MULTS_3_2(53)<=signed(MULTS_2_3(53)(PERCISION) & MULTS_2_3(53)(PERCISION downto 1))+signed(MULTS_2_4(53)(PERCISION) & MULTS_2_4(53)(PERCISION downto 1));
			MULTS_3_2(54)<=signed(MULTS_2_3(54)(PERCISION) & MULTS_2_3(54)(PERCISION downto 1))+signed(MULTS_2_4(54)(PERCISION) & MULTS_2_4(54)(PERCISION downto 1));
			MULTS_3_2(55)<=signed(MULTS_2_3(55)(PERCISION) & MULTS_2_3(55)(PERCISION downto 1))+signed(MULTS_2_4(55)(PERCISION) & MULTS_2_4(55)(PERCISION downto 1));
			MULTS_3_2(56)<=signed(MULTS_2_3(56)(PERCISION) & MULTS_2_3(56)(PERCISION downto 1))+signed(MULTS_2_4(56)(PERCISION) & MULTS_2_4(56)(PERCISION downto 1));
			MULTS_3_2(57)<=signed(MULTS_2_3(57)(PERCISION) & MULTS_2_3(57)(PERCISION downto 1))+signed(MULTS_2_4(57)(PERCISION) & MULTS_2_4(57)(PERCISION downto 1));
			MULTS_3_2(58)<=signed(MULTS_2_3(58)(PERCISION) & MULTS_2_3(58)(PERCISION downto 1))+signed(MULTS_2_4(58)(PERCISION) & MULTS_2_4(58)(PERCISION downto 1));
			MULTS_3_2(59)<=signed(MULTS_2_3(59)(PERCISION) & MULTS_2_3(59)(PERCISION downto 1))+signed(MULTS_2_4(59)(PERCISION) & MULTS_2_4(59)(PERCISION downto 1));
			MULTS_3_2(60)<=signed(MULTS_2_3(60)(PERCISION) & MULTS_2_3(60)(PERCISION downto 1))+signed(MULTS_2_4(60)(PERCISION) & MULTS_2_4(60)(PERCISION downto 1));
			MULTS_3_2(61)<=signed(MULTS_2_3(61)(PERCISION) & MULTS_2_3(61)(PERCISION downto 1))+signed(MULTS_2_4(61)(PERCISION) & MULTS_2_4(61)(PERCISION downto 1));
			MULTS_3_2(62)<=signed(MULTS_2_3(62)(PERCISION) & MULTS_2_3(62)(PERCISION downto 1))+signed(MULTS_2_4(62)(PERCISION) & MULTS_2_4(62)(PERCISION downto 1));
			MULTS_3_2(63)<=signed(MULTS_2_3(63)(PERCISION) & MULTS_2_3(63)(PERCISION downto 1))+signed(MULTS_2_4(63)(PERCISION) & MULTS_2_4(63)(PERCISION downto 1));
			MULTS_3_2(64)<=signed(MULTS_2_3(64)(PERCISION) & MULTS_2_3(64)(PERCISION downto 1))+signed(MULTS_2_4(64)(PERCISION) & MULTS_2_4(64)(PERCISION downto 1));
			MULTS_3_2(65)<=signed(MULTS_2_3(65)(PERCISION) & MULTS_2_3(65)(PERCISION downto 1))+signed(MULTS_2_4(65)(PERCISION) & MULTS_2_4(65)(PERCISION downto 1));
			MULTS_3_2(66)<=signed(MULTS_2_3(66)(PERCISION) & MULTS_2_3(66)(PERCISION downto 1))+signed(MULTS_2_4(66)(PERCISION) & MULTS_2_4(66)(PERCISION downto 1));
			MULTS_3_2(67)<=signed(MULTS_2_3(67)(PERCISION) & MULTS_2_3(67)(PERCISION downto 1))+signed(MULTS_2_4(67)(PERCISION) & MULTS_2_4(67)(PERCISION downto 1));
			MULTS_3_2(68)<=signed(MULTS_2_3(68)(PERCISION) & MULTS_2_3(68)(PERCISION downto 1))+signed(MULTS_2_4(68)(PERCISION) & MULTS_2_4(68)(PERCISION downto 1));
			MULTS_3_2(69)<=signed(MULTS_2_3(69)(PERCISION) & MULTS_2_3(69)(PERCISION downto 1))+signed(MULTS_2_4(69)(PERCISION) & MULTS_2_4(69)(PERCISION downto 1));
			MULTS_3_2(70)<=signed(MULTS_2_3(70)(PERCISION) & MULTS_2_3(70)(PERCISION downto 1))+signed(MULTS_2_4(70)(PERCISION) & MULTS_2_4(70)(PERCISION downto 1));
			MULTS_3_2(71)<=signed(MULTS_2_3(71)(PERCISION) & MULTS_2_3(71)(PERCISION downto 1))+signed(MULTS_2_4(71)(PERCISION) & MULTS_2_4(71)(PERCISION downto 1));
			MULTS_3_2(72)<=signed(MULTS_2_3(72)(PERCISION) & MULTS_2_3(72)(PERCISION downto 1))+signed(MULTS_2_4(72)(PERCISION) & MULTS_2_4(72)(PERCISION downto 1));
			MULTS_3_2(73)<=signed(MULTS_2_3(73)(PERCISION) & MULTS_2_3(73)(PERCISION downto 1))+signed(MULTS_2_4(73)(PERCISION) & MULTS_2_4(73)(PERCISION downto 1));
			MULTS_3_2(74)<=signed(MULTS_2_3(74)(PERCISION) & MULTS_2_3(74)(PERCISION downto 1))+signed(MULTS_2_4(74)(PERCISION) & MULTS_2_4(74)(PERCISION downto 1));
			MULTS_3_2(75)<=signed(MULTS_2_3(75)(PERCISION) & MULTS_2_3(75)(PERCISION downto 1))+signed(MULTS_2_4(75)(PERCISION) & MULTS_2_4(75)(PERCISION downto 1));
			MULTS_3_2(76)<=signed(MULTS_2_3(76)(PERCISION) & MULTS_2_3(76)(PERCISION downto 1))+signed(MULTS_2_4(76)(PERCISION) & MULTS_2_4(76)(PERCISION downto 1));
			MULTS_3_2(77)<=signed(MULTS_2_3(77)(PERCISION) & MULTS_2_3(77)(PERCISION downto 1))+signed(MULTS_2_4(77)(PERCISION) & MULTS_2_4(77)(PERCISION downto 1));
			MULTS_3_2(78)<=signed(MULTS_2_3(78)(PERCISION) & MULTS_2_3(78)(PERCISION downto 1))+signed(MULTS_2_4(78)(PERCISION) & MULTS_2_4(78)(PERCISION downto 1));
			MULTS_3_2(79)<=signed(MULTS_2_3(79)(PERCISION) & MULTS_2_3(79)(PERCISION downto 1))+signed(MULTS_2_4(79)(PERCISION) & MULTS_2_4(79)(PERCISION downto 1));
			MULTS_3_2(80)<=signed(MULTS_2_3(80)(PERCISION) & MULTS_2_3(80)(PERCISION downto 1))+signed(MULTS_2_4(80)(PERCISION) & MULTS_2_4(80)(PERCISION downto 1));
			MULTS_3_2(81)<=signed(MULTS_2_3(81)(PERCISION) & MULTS_2_3(81)(PERCISION downto 1))+signed(MULTS_2_4(81)(PERCISION) & MULTS_2_4(81)(PERCISION downto 1));
			MULTS_3_2(82)<=signed(MULTS_2_3(82)(PERCISION) & MULTS_2_3(82)(PERCISION downto 1))+signed(MULTS_2_4(82)(PERCISION) & MULTS_2_4(82)(PERCISION downto 1));
			MULTS_3_2(83)<=signed(MULTS_2_3(83)(PERCISION) & MULTS_2_3(83)(PERCISION downto 1))+signed(MULTS_2_4(83)(PERCISION) & MULTS_2_4(83)(PERCISION downto 1));

			MULTS_3_3(0)<=signed(MULTS_2_5(0)(PERCISION) & MULTS_2_5(0)(PERCISION downto 1))+signed(MULTS_2_6(0)(PERCISION) & MULTS_2_6(0)(PERCISION downto 1));
			MULTS_3_3(1)<=signed(MULTS_2_5(1)(PERCISION) & MULTS_2_5(1)(PERCISION downto 1))+signed(MULTS_2_6(1)(PERCISION) & MULTS_2_6(1)(PERCISION downto 1));
			MULTS_3_3(2)<=signed(MULTS_2_5(2)(PERCISION) & MULTS_2_5(2)(PERCISION downto 1))+signed(MULTS_2_6(2)(PERCISION) & MULTS_2_6(2)(PERCISION downto 1));
			MULTS_3_3(3)<=signed(MULTS_2_5(3)(PERCISION) & MULTS_2_5(3)(PERCISION downto 1))+signed(MULTS_2_6(3)(PERCISION) & MULTS_2_6(3)(PERCISION downto 1));
			MULTS_3_3(4)<=signed(MULTS_2_5(4)(PERCISION) & MULTS_2_5(4)(PERCISION downto 1))+signed(MULTS_2_6(4)(PERCISION) & MULTS_2_6(4)(PERCISION downto 1));
			MULTS_3_3(5)<=signed(MULTS_2_5(5)(PERCISION) & MULTS_2_5(5)(PERCISION downto 1))+signed(MULTS_2_6(5)(PERCISION) & MULTS_2_6(5)(PERCISION downto 1));
			MULTS_3_3(6)<=signed(MULTS_2_5(6)(PERCISION) & MULTS_2_5(6)(PERCISION downto 1))+signed(MULTS_2_6(6)(PERCISION) & MULTS_2_6(6)(PERCISION downto 1));
			MULTS_3_3(7)<=signed(MULTS_2_5(7)(PERCISION) & MULTS_2_5(7)(PERCISION downto 1))+signed(MULTS_2_6(7)(PERCISION) & MULTS_2_6(7)(PERCISION downto 1));
			MULTS_3_3(8)<=signed(MULTS_2_5(8)(PERCISION) & MULTS_2_5(8)(PERCISION downto 1))+signed(MULTS_2_6(8)(PERCISION) & MULTS_2_6(8)(PERCISION downto 1));
			MULTS_3_3(9)<=signed(MULTS_2_5(9)(PERCISION) & MULTS_2_5(9)(PERCISION downto 1))+signed(MULTS_2_6(9)(PERCISION) & MULTS_2_6(9)(PERCISION downto 1));
			MULTS_3_3(10)<=signed(MULTS_2_5(10)(PERCISION) & MULTS_2_5(10)(PERCISION downto 1))+signed(MULTS_2_6(10)(PERCISION) & MULTS_2_6(10)(PERCISION downto 1));
			MULTS_3_3(11)<=signed(MULTS_2_5(11)(PERCISION) & MULTS_2_5(11)(PERCISION downto 1))+signed(MULTS_2_6(11)(PERCISION) & MULTS_2_6(11)(PERCISION downto 1));
			MULTS_3_3(12)<=signed(MULTS_2_5(12)(PERCISION) & MULTS_2_5(12)(PERCISION downto 1))+signed(MULTS_2_6(12)(PERCISION) & MULTS_2_6(12)(PERCISION downto 1));
			MULTS_3_3(13)<=signed(MULTS_2_5(13)(PERCISION) & MULTS_2_5(13)(PERCISION downto 1))+signed(MULTS_2_6(13)(PERCISION) & MULTS_2_6(13)(PERCISION downto 1));
			MULTS_3_3(14)<=signed(MULTS_2_5(14)(PERCISION) & MULTS_2_5(14)(PERCISION downto 1))+signed(MULTS_2_6(14)(PERCISION) & MULTS_2_6(14)(PERCISION downto 1));
			MULTS_3_3(15)<=signed(MULTS_2_5(15)(PERCISION) & MULTS_2_5(15)(PERCISION downto 1))+signed(MULTS_2_6(15)(PERCISION) & MULTS_2_6(15)(PERCISION downto 1));
			MULTS_3_3(16)<=signed(MULTS_2_5(16)(PERCISION) & MULTS_2_5(16)(PERCISION downto 1))+signed(MULTS_2_6(16)(PERCISION) & MULTS_2_6(16)(PERCISION downto 1));
			MULTS_3_3(17)<=signed(MULTS_2_5(17)(PERCISION) & MULTS_2_5(17)(PERCISION downto 1))+signed(MULTS_2_6(17)(PERCISION) & MULTS_2_6(17)(PERCISION downto 1));
			MULTS_3_3(18)<=signed(MULTS_2_5(18)(PERCISION) & MULTS_2_5(18)(PERCISION downto 1))+signed(MULTS_2_6(18)(PERCISION) & MULTS_2_6(18)(PERCISION downto 1));
			MULTS_3_3(19)<=signed(MULTS_2_5(19)(PERCISION) & MULTS_2_5(19)(PERCISION downto 1))+signed(MULTS_2_6(19)(PERCISION) & MULTS_2_6(19)(PERCISION downto 1));
			MULTS_3_3(20)<=signed(MULTS_2_5(20)(PERCISION) & MULTS_2_5(20)(PERCISION downto 1))+signed(MULTS_2_6(20)(PERCISION) & MULTS_2_6(20)(PERCISION downto 1));
			MULTS_3_3(21)<=signed(MULTS_2_5(21)(PERCISION) & MULTS_2_5(21)(PERCISION downto 1))+signed(MULTS_2_6(21)(PERCISION) & MULTS_2_6(21)(PERCISION downto 1));
			MULTS_3_3(22)<=signed(MULTS_2_5(22)(PERCISION) & MULTS_2_5(22)(PERCISION downto 1))+signed(MULTS_2_6(22)(PERCISION) & MULTS_2_6(22)(PERCISION downto 1));
			MULTS_3_3(23)<=signed(MULTS_2_5(23)(PERCISION) & MULTS_2_5(23)(PERCISION downto 1))+signed(MULTS_2_6(23)(PERCISION) & MULTS_2_6(23)(PERCISION downto 1));
			MULTS_3_3(24)<=signed(MULTS_2_5(24)(PERCISION) & MULTS_2_5(24)(PERCISION downto 1))+signed(MULTS_2_6(24)(PERCISION) & MULTS_2_6(24)(PERCISION downto 1));
			MULTS_3_3(25)<=signed(MULTS_2_5(25)(PERCISION) & MULTS_2_5(25)(PERCISION downto 1))+signed(MULTS_2_6(25)(PERCISION) & MULTS_2_6(25)(PERCISION downto 1));
			MULTS_3_3(26)<=signed(MULTS_2_5(26)(PERCISION) & MULTS_2_5(26)(PERCISION downto 1))+signed(MULTS_2_6(26)(PERCISION) & MULTS_2_6(26)(PERCISION downto 1));
			MULTS_3_3(27)<=signed(MULTS_2_5(27)(PERCISION) & MULTS_2_5(27)(PERCISION downto 1))+signed(MULTS_2_6(27)(PERCISION) & MULTS_2_6(27)(PERCISION downto 1));
			MULTS_3_3(28)<=signed(MULTS_2_5(28)(PERCISION) & MULTS_2_5(28)(PERCISION downto 1))+signed(MULTS_2_6(28)(PERCISION) & MULTS_2_6(28)(PERCISION downto 1));
			MULTS_3_3(29)<=signed(MULTS_2_5(29)(PERCISION) & MULTS_2_5(29)(PERCISION downto 1))+signed(MULTS_2_6(29)(PERCISION) & MULTS_2_6(29)(PERCISION downto 1));
			MULTS_3_3(30)<=signed(MULTS_2_5(30)(PERCISION) & MULTS_2_5(30)(PERCISION downto 1))+signed(MULTS_2_6(30)(PERCISION) & MULTS_2_6(30)(PERCISION downto 1));
			MULTS_3_3(31)<=signed(MULTS_2_5(31)(PERCISION) & MULTS_2_5(31)(PERCISION downto 1))+signed(MULTS_2_6(31)(PERCISION) & MULTS_2_6(31)(PERCISION downto 1));
			MULTS_3_3(32)<=signed(MULTS_2_5(32)(PERCISION) & MULTS_2_5(32)(PERCISION downto 1))+signed(MULTS_2_6(32)(PERCISION) & MULTS_2_6(32)(PERCISION downto 1));
			MULTS_3_3(33)<=signed(MULTS_2_5(33)(PERCISION) & MULTS_2_5(33)(PERCISION downto 1))+signed(MULTS_2_6(33)(PERCISION) & MULTS_2_6(33)(PERCISION downto 1));
			MULTS_3_3(34)<=signed(MULTS_2_5(34)(PERCISION) & MULTS_2_5(34)(PERCISION downto 1))+signed(MULTS_2_6(34)(PERCISION) & MULTS_2_6(34)(PERCISION downto 1));
			MULTS_3_3(35)<=signed(MULTS_2_5(35)(PERCISION) & MULTS_2_5(35)(PERCISION downto 1))+signed(MULTS_2_6(35)(PERCISION) & MULTS_2_6(35)(PERCISION downto 1));
			MULTS_3_3(36)<=signed(MULTS_2_5(36)(PERCISION) & MULTS_2_5(36)(PERCISION downto 1))+signed(MULTS_2_6(36)(PERCISION) & MULTS_2_6(36)(PERCISION downto 1));
			MULTS_3_3(37)<=signed(MULTS_2_5(37)(PERCISION) & MULTS_2_5(37)(PERCISION downto 1))+signed(MULTS_2_6(37)(PERCISION) & MULTS_2_6(37)(PERCISION downto 1));
			MULTS_3_3(38)<=signed(MULTS_2_5(38)(PERCISION) & MULTS_2_5(38)(PERCISION downto 1))+signed(MULTS_2_6(38)(PERCISION) & MULTS_2_6(38)(PERCISION downto 1));
			MULTS_3_3(39)<=signed(MULTS_2_5(39)(PERCISION) & MULTS_2_5(39)(PERCISION downto 1))+signed(MULTS_2_6(39)(PERCISION) & MULTS_2_6(39)(PERCISION downto 1));
			MULTS_3_3(40)<=signed(MULTS_2_5(40)(PERCISION) & MULTS_2_5(40)(PERCISION downto 1))+signed(MULTS_2_6(40)(PERCISION) & MULTS_2_6(40)(PERCISION downto 1));
			MULTS_3_3(41)<=signed(MULTS_2_5(41)(PERCISION) & MULTS_2_5(41)(PERCISION downto 1))+signed(MULTS_2_6(41)(PERCISION) & MULTS_2_6(41)(PERCISION downto 1));
			MULTS_3_3(42)<=signed(MULTS_2_5(42)(PERCISION) & MULTS_2_5(42)(PERCISION downto 1))+signed(MULTS_2_6(42)(PERCISION) & MULTS_2_6(42)(PERCISION downto 1));
			MULTS_3_3(43)<=signed(MULTS_2_5(43)(PERCISION) & MULTS_2_5(43)(PERCISION downto 1))+signed(MULTS_2_6(43)(PERCISION) & MULTS_2_6(43)(PERCISION downto 1));
			MULTS_3_3(44)<=signed(MULTS_2_5(44)(PERCISION) & MULTS_2_5(44)(PERCISION downto 1))+signed(MULTS_2_6(44)(PERCISION) & MULTS_2_6(44)(PERCISION downto 1));
			MULTS_3_3(45)<=signed(MULTS_2_5(45)(PERCISION) & MULTS_2_5(45)(PERCISION downto 1))+signed(MULTS_2_6(45)(PERCISION) & MULTS_2_6(45)(PERCISION downto 1));
			MULTS_3_3(46)<=signed(MULTS_2_5(46)(PERCISION) & MULTS_2_5(46)(PERCISION downto 1))+signed(MULTS_2_6(46)(PERCISION) & MULTS_2_6(46)(PERCISION downto 1));
			MULTS_3_3(47)<=signed(MULTS_2_5(47)(PERCISION) & MULTS_2_5(47)(PERCISION downto 1))+signed(MULTS_2_6(47)(PERCISION) & MULTS_2_6(47)(PERCISION downto 1));
			MULTS_3_3(48)<=signed(MULTS_2_5(48)(PERCISION) & MULTS_2_5(48)(PERCISION downto 1))+signed(MULTS_2_6(48)(PERCISION) & MULTS_2_6(48)(PERCISION downto 1));
			MULTS_3_3(49)<=signed(MULTS_2_5(49)(PERCISION) & MULTS_2_5(49)(PERCISION downto 1))+signed(MULTS_2_6(49)(PERCISION) & MULTS_2_6(49)(PERCISION downto 1));
			MULTS_3_3(50)<=signed(MULTS_2_5(50)(PERCISION) & MULTS_2_5(50)(PERCISION downto 1))+signed(MULTS_2_6(50)(PERCISION) & MULTS_2_6(50)(PERCISION downto 1));
			MULTS_3_3(51)<=signed(MULTS_2_5(51)(PERCISION) & MULTS_2_5(51)(PERCISION downto 1))+signed(MULTS_2_6(51)(PERCISION) & MULTS_2_6(51)(PERCISION downto 1));
			MULTS_3_3(52)<=signed(MULTS_2_5(52)(PERCISION) & MULTS_2_5(52)(PERCISION downto 1))+signed(MULTS_2_6(52)(PERCISION) & MULTS_2_6(52)(PERCISION downto 1));
			MULTS_3_3(53)<=signed(MULTS_2_5(53)(PERCISION) & MULTS_2_5(53)(PERCISION downto 1))+signed(MULTS_2_6(53)(PERCISION) & MULTS_2_6(53)(PERCISION downto 1));
			MULTS_3_3(54)<=signed(MULTS_2_5(54)(PERCISION) & MULTS_2_5(54)(PERCISION downto 1))+signed(MULTS_2_6(54)(PERCISION) & MULTS_2_6(54)(PERCISION downto 1));
			MULTS_3_3(55)<=signed(MULTS_2_5(55)(PERCISION) & MULTS_2_5(55)(PERCISION downto 1))+signed(MULTS_2_6(55)(PERCISION) & MULTS_2_6(55)(PERCISION downto 1));
			MULTS_3_3(56)<=signed(MULTS_2_5(56)(PERCISION) & MULTS_2_5(56)(PERCISION downto 1))+signed(MULTS_2_6(56)(PERCISION) & MULTS_2_6(56)(PERCISION downto 1));
			MULTS_3_3(57)<=signed(MULTS_2_5(57)(PERCISION) & MULTS_2_5(57)(PERCISION downto 1))+signed(MULTS_2_6(57)(PERCISION) & MULTS_2_6(57)(PERCISION downto 1));
			MULTS_3_3(58)<=signed(MULTS_2_5(58)(PERCISION) & MULTS_2_5(58)(PERCISION downto 1))+signed(MULTS_2_6(58)(PERCISION) & MULTS_2_6(58)(PERCISION downto 1));
			MULTS_3_3(59)<=signed(MULTS_2_5(59)(PERCISION) & MULTS_2_5(59)(PERCISION downto 1))+signed(MULTS_2_6(59)(PERCISION) & MULTS_2_6(59)(PERCISION downto 1));
			MULTS_3_3(60)<=signed(MULTS_2_5(60)(PERCISION) & MULTS_2_5(60)(PERCISION downto 1))+signed(MULTS_2_6(60)(PERCISION) & MULTS_2_6(60)(PERCISION downto 1));
			MULTS_3_3(61)<=signed(MULTS_2_5(61)(PERCISION) & MULTS_2_5(61)(PERCISION downto 1))+signed(MULTS_2_6(61)(PERCISION) & MULTS_2_6(61)(PERCISION downto 1));
			MULTS_3_3(62)<=signed(MULTS_2_5(62)(PERCISION) & MULTS_2_5(62)(PERCISION downto 1))+signed(MULTS_2_6(62)(PERCISION) & MULTS_2_6(62)(PERCISION downto 1));
			MULTS_3_3(63)<=signed(MULTS_2_5(63)(PERCISION) & MULTS_2_5(63)(PERCISION downto 1))+signed(MULTS_2_6(63)(PERCISION) & MULTS_2_6(63)(PERCISION downto 1));
			MULTS_3_3(64)<=signed(MULTS_2_5(64)(PERCISION) & MULTS_2_5(64)(PERCISION downto 1))+signed(MULTS_2_6(64)(PERCISION) & MULTS_2_6(64)(PERCISION downto 1));
			MULTS_3_3(65)<=signed(MULTS_2_5(65)(PERCISION) & MULTS_2_5(65)(PERCISION downto 1))+signed(MULTS_2_6(65)(PERCISION) & MULTS_2_6(65)(PERCISION downto 1));
			MULTS_3_3(66)<=signed(MULTS_2_5(66)(PERCISION) & MULTS_2_5(66)(PERCISION downto 1))+signed(MULTS_2_6(66)(PERCISION) & MULTS_2_6(66)(PERCISION downto 1));
			MULTS_3_3(67)<=signed(MULTS_2_5(67)(PERCISION) & MULTS_2_5(67)(PERCISION downto 1))+signed(MULTS_2_6(67)(PERCISION) & MULTS_2_6(67)(PERCISION downto 1));
			MULTS_3_3(68)<=signed(MULTS_2_5(68)(PERCISION) & MULTS_2_5(68)(PERCISION downto 1))+signed(MULTS_2_6(68)(PERCISION) & MULTS_2_6(68)(PERCISION downto 1));
			MULTS_3_3(69)<=signed(MULTS_2_5(69)(PERCISION) & MULTS_2_5(69)(PERCISION downto 1))+signed(MULTS_2_6(69)(PERCISION) & MULTS_2_6(69)(PERCISION downto 1));
			MULTS_3_3(70)<=signed(MULTS_2_5(70)(PERCISION) & MULTS_2_5(70)(PERCISION downto 1))+signed(MULTS_2_6(70)(PERCISION) & MULTS_2_6(70)(PERCISION downto 1));
			MULTS_3_3(71)<=signed(MULTS_2_5(71)(PERCISION) & MULTS_2_5(71)(PERCISION downto 1))+signed(MULTS_2_6(71)(PERCISION) & MULTS_2_6(71)(PERCISION downto 1));
			MULTS_3_3(72)<=signed(MULTS_2_5(72)(PERCISION) & MULTS_2_5(72)(PERCISION downto 1))+signed(MULTS_2_6(72)(PERCISION) & MULTS_2_6(72)(PERCISION downto 1));
			MULTS_3_3(73)<=signed(MULTS_2_5(73)(PERCISION) & MULTS_2_5(73)(PERCISION downto 1))+signed(MULTS_2_6(73)(PERCISION) & MULTS_2_6(73)(PERCISION downto 1));
			MULTS_3_3(74)<=signed(MULTS_2_5(74)(PERCISION) & MULTS_2_5(74)(PERCISION downto 1))+signed(MULTS_2_6(74)(PERCISION) & MULTS_2_6(74)(PERCISION downto 1));
			MULTS_3_3(75)<=signed(MULTS_2_5(75)(PERCISION) & MULTS_2_5(75)(PERCISION downto 1))+signed(MULTS_2_6(75)(PERCISION) & MULTS_2_6(75)(PERCISION downto 1));
			MULTS_3_3(76)<=signed(MULTS_2_5(76)(PERCISION) & MULTS_2_5(76)(PERCISION downto 1))+signed(MULTS_2_6(76)(PERCISION) & MULTS_2_6(76)(PERCISION downto 1));
			MULTS_3_3(77)<=signed(MULTS_2_5(77)(PERCISION) & MULTS_2_5(77)(PERCISION downto 1))+signed(MULTS_2_6(77)(PERCISION) & MULTS_2_6(77)(PERCISION downto 1));
			MULTS_3_3(78)<=signed(MULTS_2_5(78)(PERCISION) & MULTS_2_5(78)(PERCISION downto 1))+signed(MULTS_2_6(78)(PERCISION) & MULTS_2_6(78)(PERCISION downto 1));
			MULTS_3_3(79)<=signed(MULTS_2_5(79)(PERCISION) & MULTS_2_5(79)(PERCISION downto 1))+signed(MULTS_2_6(79)(PERCISION) & MULTS_2_6(79)(PERCISION downto 1));
			MULTS_3_3(80)<=signed(MULTS_2_5(80)(PERCISION) & MULTS_2_5(80)(PERCISION downto 1))+signed(MULTS_2_6(80)(PERCISION) & MULTS_2_6(80)(PERCISION downto 1));
			MULTS_3_3(81)<=signed(MULTS_2_5(81)(PERCISION) & MULTS_2_5(81)(PERCISION downto 1))+signed(MULTS_2_6(81)(PERCISION) & MULTS_2_6(81)(PERCISION downto 1));
			MULTS_3_3(82)<=signed(MULTS_2_5(82)(PERCISION) & MULTS_2_5(82)(PERCISION downto 1))+signed(MULTS_2_6(82)(PERCISION) & MULTS_2_6(82)(PERCISION downto 1));
			MULTS_3_3(83)<=signed(MULTS_2_5(83)(PERCISION) & MULTS_2_5(83)(PERCISION downto 1))+signed(MULTS_2_6(83)(PERCISION) & MULTS_2_6(83)(PERCISION downto 1));

			MULTS_3_4(0)<=signed(MULTS_2_7(0)(PERCISION) & MULTS_2_7(0)(PERCISION downto 1))+signed(MULTS_2_8(0)(PERCISION) & MULTS_2_8(0)(PERCISION downto 1));
			MULTS_3_4(1)<=signed(MULTS_2_7(1)(PERCISION) & MULTS_2_7(1)(PERCISION downto 1))+signed(MULTS_2_8(1)(PERCISION) & MULTS_2_8(1)(PERCISION downto 1));
			MULTS_3_4(2)<=signed(MULTS_2_7(2)(PERCISION) & MULTS_2_7(2)(PERCISION downto 1))+signed(MULTS_2_8(2)(PERCISION) & MULTS_2_8(2)(PERCISION downto 1));
			MULTS_3_4(3)<=signed(MULTS_2_7(3)(PERCISION) & MULTS_2_7(3)(PERCISION downto 1))+signed(MULTS_2_8(3)(PERCISION) & MULTS_2_8(3)(PERCISION downto 1));
			MULTS_3_4(4)<=signed(MULTS_2_7(4)(PERCISION) & MULTS_2_7(4)(PERCISION downto 1))+signed(MULTS_2_8(4)(PERCISION) & MULTS_2_8(4)(PERCISION downto 1));
			MULTS_3_4(5)<=signed(MULTS_2_7(5)(PERCISION) & MULTS_2_7(5)(PERCISION downto 1))+signed(MULTS_2_8(5)(PERCISION) & MULTS_2_8(5)(PERCISION downto 1));
			MULTS_3_4(6)<=signed(MULTS_2_7(6)(PERCISION) & MULTS_2_7(6)(PERCISION downto 1))+signed(MULTS_2_8(6)(PERCISION) & MULTS_2_8(6)(PERCISION downto 1));
			MULTS_3_4(7)<=signed(MULTS_2_7(7)(PERCISION) & MULTS_2_7(7)(PERCISION downto 1))+signed(MULTS_2_8(7)(PERCISION) & MULTS_2_8(7)(PERCISION downto 1));
			MULTS_3_4(8)<=signed(MULTS_2_7(8)(PERCISION) & MULTS_2_7(8)(PERCISION downto 1))+signed(MULTS_2_8(8)(PERCISION) & MULTS_2_8(8)(PERCISION downto 1));
			MULTS_3_4(9)<=signed(MULTS_2_7(9)(PERCISION) & MULTS_2_7(9)(PERCISION downto 1))+signed(MULTS_2_8(9)(PERCISION) & MULTS_2_8(9)(PERCISION downto 1));
			MULTS_3_4(10)<=signed(MULTS_2_7(10)(PERCISION) & MULTS_2_7(10)(PERCISION downto 1))+signed(MULTS_2_8(10)(PERCISION) & MULTS_2_8(10)(PERCISION downto 1));
			MULTS_3_4(11)<=signed(MULTS_2_7(11)(PERCISION) & MULTS_2_7(11)(PERCISION downto 1))+signed(MULTS_2_8(11)(PERCISION) & MULTS_2_8(11)(PERCISION downto 1));
			MULTS_3_4(12)<=signed(MULTS_2_7(12)(PERCISION) & MULTS_2_7(12)(PERCISION downto 1))+signed(MULTS_2_8(12)(PERCISION) & MULTS_2_8(12)(PERCISION downto 1));
			MULTS_3_4(13)<=signed(MULTS_2_7(13)(PERCISION) & MULTS_2_7(13)(PERCISION downto 1))+signed(MULTS_2_8(13)(PERCISION) & MULTS_2_8(13)(PERCISION downto 1));
			MULTS_3_4(14)<=signed(MULTS_2_7(14)(PERCISION) & MULTS_2_7(14)(PERCISION downto 1))+signed(MULTS_2_8(14)(PERCISION) & MULTS_2_8(14)(PERCISION downto 1));
			MULTS_3_4(15)<=signed(MULTS_2_7(15)(PERCISION) & MULTS_2_7(15)(PERCISION downto 1))+signed(MULTS_2_8(15)(PERCISION) & MULTS_2_8(15)(PERCISION downto 1));
			MULTS_3_4(16)<=signed(MULTS_2_7(16)(PERCISION) & MULTS_2_7(16)(PERCISION downto 1))+signed(MULTS_2_8(16)(PERCISION) & MULTS_2_8(16)(PERCISION downto 1));
			MULTS_3_4(17)<=signed(MULTS_2_7(17)(PERCISION) & MULTS_2_7(17)(PERCISION downto 1))+signed(MULTS_2_8(17)(PERCISION) & MULTS_2_8(17)(PERCISION downto 1));
			MULTS_3_4(18)<=signed(MULTS_2_7(18)(PERCISION) & MULTS_2_7(18)(PERCISION downto 1))+signed(MULTS_2_8(18)(PERCISION) & MULTS_2_8(18)(PERCISION downto 1));
			MULTS_3_4(19)<=signed(MULTS_2_7(19)(PERCISION) & MULTS_2_7(19)(PERCISION downto 1))+signed(MULTS_2_8(19)(PERCISION) & MULTS_2_8(19)(PERCISION downto 1));
			MULTS_3_4(20)<=signed(MULTS_2_7(20)(PERCISION) & MULTS_2_7(20)(PERCISION downto 1))+signed(MULTS_2_8(20)(PERCISION) & MULTS_2_8(20)(PERCISION downto 1));
			MULTS_3_4(21)<=signed(MULTS_2_7(21)(PERCISION) & MULTS_2_7(21)(PERCISION downto 1))+signed(MULTS_2_8(21)(PERCISION) & MULTS_2_8(21)(PERCISION downto 1));
			MULTS_3_4(22)<=signed(MULTS_2_7(22)(PERCISION) & MULTS_2_7(22)(PERCISION downto 1))+signed(MULTS_2_8(22)(PERCISION) & MULTS_2_8(22)(PERCISION downto 1));
			MULTS_3_4(23)<=signed(MULTS_2_7(23)(PERCISION) & MULTS_2_7(23)(PERCISION downto 1))+signed(MULTS_2_8(23)(PERCISION) & MULTS_2_8(23)(PERCISION downto 1));
			MULTS_3_4(24)<=signed(MULTS_2_7(24)(PERCISION) & MULTS_2_7(24)(PERCISION downto 1))+signed(MULTS_2_8(24)(PERCISION) & MULTS_2_8(24)(PERCISION downto 1));
			MULTS_3_4(25)<=signed(MULTS_2_7(25)(PERCISION) & MULTS_2_7(25)(PERCISION downto 1))+signed(MULTS_2_8(25)(PERCISION) & MULTS_2_8(25)(PERCISION downto 1));
			MULTS_3_4(26)<=signed(MULTS_2_7(26)(PERCISION) & MULTS_2_7(26)(PERCISION downto 1))+signed(MULTS_2_8(26)(PERCISION) & MULTS_2_8(26)(PERCISION downto 1));
			MULTS_3_4(27)<=signed(MULTS_2_7(27)(PERCISION) & MULTS_2_7(27)(PERCISION downto 1))+signed(MULTS_2_8(27)(PERCISION) & MULTS_2_8(27)(PERCISION downto 1));
			MULTS_3_4(28)<=signed(MULTS_2_7(28)(PERCISION) & MULTS_2_7(28)(PERCISION downto 1))+signed(MULTS_2_8(28)(PERCISION) & MULTS_2_8(28)(PERCISION downto 1));
			MULTS_3_4(29)<=signed(MULTS_2_7(29)(PERCISION) & MULTS_2_7(29)(PERCISION downto 1))+signed(MULTS_2_8(29)(PERCISION) & MULTS_2_8(29)(PERCISION downto 1));
			MULTS_3_4(30)<=signed(MULTS_2_7(30)(PERCISION) & MULTS_2_7(30)(PERCISION downto 1))+signed(MULTS_2_8(30)(PERCISION) & MULTS_2_8(30)(PERCISION downto 1));
			MULTS_3_4(31)<=signed(MULTS_2_7(31)(PERCISION) & MULTS_2_7(31)(PERCISION downto 1))+signed(MULTS_2_8(31)(PERCISION) & MULTS_2_8(31)(PERCISION downto 1));
			MULTS_3_4(32)<=signed(MULTS_2_7(32)(PERCISION) & MULTS_2_7(32)(PERCISION downto 1))+signed(MULTS_2_8(32)(PERCISION) & MULTS_2_8(32)(PERCISION downto 1));
			MULTS_3_4(33)<=signed(MULTS_2_7(33)(PERCISION) & MULTS_2_7(33)(PERCISION downto 1))+signed(MULTS_2_8(33)(PERCISION) & MULTS_2_8(33)(PERCISION downto 1));
			MULTS_3_4(34)<=signed(MULTS_2_7(34)(PERCISION) & MULTS_2_7(34)(PERCISION downto 1))+signed(MULTS_2_8(34)(PERCISION) & MULTS_2_8(34)(PERCISION downto 1));
			MULTS_3_4(35)<=signed(MULTS_2_7(35)(PERCISION) & MULTS_2_7(35)(PERCISION downto 1))+signed(MULTS_2_8(35)(PERCISION) & MULTS_2_8(35)(PERCISION downto 1));
			MULTS_3_4(36)<=signed(MULTS_2_7(36)(PERCISION) & MULTS_2_7(36)(PERCISION downto 1))+signed(MULTS_2_8(36)(PERCISION) & MULTS_2_8(36)(PERCISION downto 1));
			MULTS_3_4(37)<=signed(MULTS_2_7(37)(PERCISION) & MULTS_2_7(37)(PERCISION downto 1))+signed(MULTS_2_8(37)(PERCISION) & MULTS_2_8(37)(PERCISION downto 1));
			MULTS_3_4(38)<=signed(MULTS_2_7(38)(PERCISION) & MULTS_2_7(38)(PERCISION downto 1))+signed(MULTS_2_8(38)(PERCISION) & MULTS_2_8(38)(PERCISION downto 1));
			MULTS_3_4(39)<=signed(MULTS_2_7(39)(PERCISION) & MULTS_2_7(39)(PERCISION downto 1))+signed(MULTS_2_8(39)(PERCISION) & MULTS_2_8(39)(PERCISION downto 1));
			MULTS_3_4(40)<=signed(MULTS_2_7(40)(PERCISION) & MULTS_2_7(40)(PERCISION downto 1))+signed(MULTS_2_8(40)(PERCISION) & MULTS_2_8(40)(PERCISION downto 1));
			MULTS_3_4(41)<=signed(MULTS_2_7(41)(PERCISION) & MULTS_2_7(41)(PERCISION downto 1))+signed(MULTS_2_8(41)(PERCISION) & MULTS_2_8(41)(PERCISION downto 1));
			MULTS_3_4(42)<=signed(MULTS_2_7(42)(PERCISION) & MULTS_2_7(42)(PERCISION downto 1))+signed(MULTS_2_8(42)(PERCISION) & MULTS_2_8(42)(PERCISION downto 1));
			MULTS_3_4(43)<=signed(MULTS_2_7(43)(PERCISION) & MULTS_2_7(43)(PERCISION downto 1))+signed(MULTS_2_8(43)(PERCISION) & MULTS_2_8(43)(PERCISION downto 1));
			MULTS_3_4(44)<=signed(MULTS_2_7(44)(PERCISION) & MULTS_2_7(44)(PERCISION downto 1))+signed(MULTS_2_8(44)(PERCISION) & MULTS_2_8(44)(PERCISION downto 1));
			MULTS_3_4(45)<=signed(MULTS_2_7(45)(PERCISION) & MULTS_2_7(45)(PERCISION downto 1))+signed(MULTS_2_8(45)(PERCISION) & MULTS_2_8(45)(PERCISION downto 1));
			MULTS_3_4(46)<=signed(MULTS_2_7(46)(PERCISION) & MULTS_2_7(46)(PERCISION downto 1))+signed(MULTS_2_8(46)(PERCISION) & MULTS_2_8(46)(PERCISION downto 1));
			MULTS_3_4(47)<=signed(MULTS_2_7(47)(PERCISION) & MULTS_2_7(47)(PERCISION downto 1))+signed(MULTS_2_8(47)(PERCISION) & MULTS_2_8(47)(PERCISION downto 1));
			MULTS_3_4(48)<=signed(MULTS_2_7(48)(PERCISION) & MULTS_2_7(48)(PERCISION downto 1))+signed(MULTS_2_8(48)(PERCISION) & MULTS_2_8(48)(PERCISION downto 1));
			MULTS_3_4(49)<=signed(MULTS_2_7(49)(PERCISION) & MULTS_2_7(49)(PERCISION downto 1))+signed(MULTS_2_8(49)(PERCISION) & MULTS_2_8(49)(PERCISION downto 1));
			MULTS_3_4(50)<=signed(MULTS_2_7(50)(PERCISION) & MULTS_2_7(50)(PERCISION downto 1))+signed(MULTS_2_8(50)(PERCISION) & MULTS_2_8(50)(PERCISION downto 1));
			MULTS_3_4(51)<=signed(MULTS_2_7(51)(PERCISION) & MULTS_2_7(51)(PERCISION downto 1))+signed(MULTS_2_8(51)(PERCISION) & MULTS_2_8(51)(PERCISION downto 1));
			MULTS_3_4(52)<=signed(MULTS_2_7(52)(PERCISION) & MULTS_2_7(52)(PERCISION downto 1))+signed(MULTS_2_8(52)(PERCISION) & MULTS_2_8(52)(PERCISION downto 1));
			MULTS_3_4(53)<=signed(MULTS_2_7(53)(PERCISION) & MULTS_2_7(53)(PERCISION downto 1))+signed(MULTS_2_8(53)(PERCISION) & MULTS_2_8(53)(PERCISION downto 1));
			MULTS_3_4(54)<=signed(MULTS_2_7(54)(PERCISION) & MULTS_2_7(54)(PERCISION downto 1))+signed(MULTS_2_8(54)(PERCISION) & MULTS_2_8(54)(PERCISION downto 1));
			MULTS_3_4(55)<=signed(MULTS_2_7(55)(PERCISION) & MULTS_2_7(55)(PERCISION downto 1))+signed(MULTS_2_8(55)(PERCISION) & MULTS_2_8(55)(PERCISION downto 1));
			MULTS_3_4(56)<=signed(MULTS_2_7(56)(PERCISION) & MULTS_2_7(56)(PERCISION downto 1))+signed(MULTS_2_8(56)(PERCISION) & MULTS_2_8(56)(PERCISION downto 1));
			MULTS_3_4(57)<=signed(MULTS_2_7(57)(PERCISION) & MULTS_2_7(57)(PERCISION downto 1))+signed(MULTS_2_8(57)(PERCISION) & MULTS_2_8(57)(PERCISION downto 1));
			MULTS_3_4(58)<=signed(MULTS_2_7(58)(PERCISION) & MULTS_2_7(58)(PERCISION downto 1))+signed(MULTS_2_8(58)(PERCISION) & MULTS_2_8(58)(PERCISION downto 1));
			MULTS_3_4(59)<=signed(MULTS_2_7(59)(PERCISION) & MULTS_2_7(59)(PERCISION downto 1))+signed(MULTS_2_8(59)(PERCISION) & MULTS_2_8(59)(PERCISION downto 1));
			MULTS_3_4(60)<=signed(MULTS_2_7(60)(PERCISION) & MULTS_2_7(60)(PERCISION downto 1))+signed(MULTS_2_8(60)(PERCISION) & MULTS_2_8(60)(PERCISION downto 1));
			MULTS_3_4(61)<=signed(MULTS_2_7(61)(PERCISION) & MULTS_2_7(61)(PERCISION downto 1))+signed(MULTS_2_8(61)(PERCISION) & MULTS_2_8(61)(PERCISION downto 1));
			MULTS_3_4(62)<=signed(MULTS_2_7(62)(PERCISION) & MULTS_2_7(62)(PERCISION downto 1))+signed(MULTS_2_8(62)(PERCISION) & MULTS_2_8(62)(PERCISION downto 1));
			MULTS_3_4(63)<=signed(MULTS_2_7(63)(PERCISION) & MULTS_2_7(63)(PERCISION downto 1))+signed(MULTS_2_8(63)(PERCISION) & MULTS_2_8(63)(PERCISION downto 1));
			MULTS_3_4(64)<=signed(MULTS_2_7(64)(PERCISION) & MULTS_2_7(64)(PERCISION downto 1))+signed(MULTS_2_8(64)(PERCISION) & MULTS_2_8(64)(PERCISION downto 1));
			MULTS_3_4(65)<=signed(MULTS_2_7(65)(PERCISION) & MULTS_2_7(65)(PERCISION downto 1))+signed(MULTS_2_8(65)(PERCISION) & MULTS_2_8(65)(PERCISION downto 1));
			MULTS_3_4(66)<=signed(MULTS_2_7(66)(PERCISION) & MULTS_2_7(66)(PERCISION downto 1))+signed(MULTS_2_8(66)(PERCISION) & MULTS_2_8(66)(PERCISION downto 1));
			MULTS_3_4(67)<=signed(MULTS_2_7(67)(PERCISION) & MULTS_2_7(67)(PERCISION downto 1))+signed(MULTS_2_8(67)(PERCISION) & MULTS_2_8(67)(PERCISION downto 1));
			MULTS_3_4(68)<=signed(MULTS_2_7(68)(PERCISION) & MULTS_2_7(68)(PERCISION downto 1))+signed(MULTS_2_8(68)(PERCISION) & MULTS_2_8(68)(PERCISION downto 1));
			MULTS_3_4(69)<=signed(MULTS_2_7(69)(PERCISION) & MULTS_2_7(69)(PERCISION downto 1))+signed(MULTS_2_8(69)(PERCISION) & MULTS_2_8(69)(PERCISION downto 1));
			MULTS_3_4(70)<=signed(MULTS_2_7(70)(PERCISION) & MULTS_2_7(70)(PERCISION downto 1))+signed(MULTS_2_8(70)(PERCISION) & MULTS_2_8(70)(PERCISION downto 1));
			MULTS_3_4(71)<=signed(MULTS_2_7(71)(PERCISION) & MULTS_2_7(71)(PERCISION downto 1))+signed(MULTS_2_8(71)(PERCISION) & MULTS_2_8(71)(PERCISION downto 1));
			MULTS_3_4(72)<=signed(MULTS_2_7(72)(PERCISION) & MULTS_2_7(72)(PERCISION downto 1))+signed(MULTS_2_8(72)(PERCISION) & MULTS_2_8(72)(PERCISION downto 1));
			MULTS_3_4(73)<=signed(MULTS_2_7(73)(PERCISION) & MULTS_2_7(73)(PERCISION downto 1))+signed(MULTS_2_8(73)(PERCISION) & MULTS_2_8(73)(PERCISION downto 1));
			MULTS_3_4(74)<=signed(MULTS_2_7(74)(PERCISION) & MULTS_2_7(74)(PERCISION downto 1))+signed(MULTS_2_8(74)(PERCISION) & MULTS_2_8(74)(PERCISION downto 1));
			MULTS_3_4(75)<=signed(MULTS_2_7(75)(PERCISION) & MULTS_2_7(75)(PERCISION downto 1))+signed(MULTS_2_8(75)(PERCISION) & MULTS_2_8(75)(PERCISION downto 1));
			MULTS_3_4(76)<=signed(MULTS_2_7(76)(PERCISION) & MULTS_2_7(76)(PERCISION downto 1))+signed(MULTS_2_8(76)(PERCISION) & MULTS_2_8(76)(PERCISION downto 1));
			MULTS_3_4(77)<=signed(MULTS_2_7(77)(PERCISION) & MULTS_2_7(77)(PERCISION downto 1))+signed(MULTS_2_8(77)(PERCISION) & MULTS_2_8(77)(PERCISION downto 1));
			MULTS_3_4(78)<=signed(MULTS_2_7(78)(PERCISION) & MULTS_2_7(78)(PERCISION downto 1))+signed(MULTS_2_8(78)(PERCISION) & MULTS_2_8(78)(PERCISION downto 1));
			MULTS_3_4(79)<=signed(MULTS_2_7(79)(PERCISION) & MULTS_2_7(79)(PERCISION downto 1))+signed(MULTS_2_8(79)(PERCISION) & MULTS_2_8(79)(PERCISION downto 1));
			MULTS_3_4(80)<=signed(MULTS_2_7(80)(PERCISION) & MULTS_2_7(80)(PERCISION downto 1))+signed(MULTS_2_8(80)(PERCISION) & MULTS_2_8(80)(PERCISION downto 1));
			MULTS_3_4(81)<=signed(MULTS_2_7(81)(PERCISION) & MULTS_2_7(81)(PERCISION downto 1))+signed(MULTS_2_8(81)(PERCISION) & MULTS_2_8(81)(PERCISION downto 1));
			MULTS_3_4(82)<=signed(MULTS_2_7(82)(PERCISION) & MULTS_2_7(82)(PERCISION downto 1))+signed(MULTS_2_8(82)(PERCISION) & MULTS_2_8(82)(PERCISION downto 1));
			MULTS_3_4(83)<=signed(MULTS_2_7(83)(PERCISION) & MULTS_2_7(83)(PERCISION downto 1))+signed(MULTS_2_8(83)(PERCISION) & MULTS_2_8(83)(PERCISION downto 1));

			MULTS_3_5(0)<=signed(MULTS_2_9(0)(PERCISION) & MULTS_2_9(0)(PERCISION downto 1))+signed(MULTS_2_10(0)(PERCISION) & MULTS_2_10(0)(PERCISION downto 1));
			MULTS_3_5(1)<=signed(MULTS_2_9(1)(PERCISION) & MULTS_2_9(1)(PERCISION downto 1))+signed(MULTS_2_10(1)(PERCISION) & MULTS_2_10(1)(PERCISION downto 1));
			MULTS_3_5(2)<=signed(MULTS_2_9(2)(PERCISION) & MULTS_2_9(2)(PERCISION downto 1))+signed(MULTS_2_10(2)(PERCISION) & MULTS_2_10(2)(PERCISION downto 1));
			MULTS_3_5(3)<=signed(MULTS_2_9(3)(PERCISION) & MULTS_2_9(3)(PERCISION downto 1))+signed(MULTS_2_10(3)(PERCISION) & MULTS_2_10(3)(PERCISION downto 1));
			MULTS_3_5(4)<=signed(MULTS_2_9(4)(PERCISION) & MULTS_2_9(4)(PERCISION downto 1))+signed(MULTS_2_10(4)(PERCISION) & MULTS_2_10(4)(PERCISION downto 1));
			MULTS_3_5(5)<=signed(MULTS_2_9(5)(PERCISION) & MULTS_2_9(5)(PERCISION downto 1))+signed(MULTS_2_10(5)(PERCISION) & MULTS_2_10(5)(PERCISION downto 1));
			MULTS_3_5(6)<=signed(MULTS_2_9(6)(PERCISION) & MULTS_2_9(6)(PERCISION downto 1))+signed(MULTS_2_10(6)(PERCISION) & MULTS_2_10(6)(PERCISION downto 1));
			MULTS_3_5(7)<=signed(MULTS_2_9(7)(PERCISION) & MULTS_2_9(7)(PERCISION downto 1))+signed(MULTS_2_10(7)(PERCISION) & MULTS_2_10(7)(PERCISION downto 1));
			MULTS_3_5(8)<=signed(MULTS_2_9(8)(PERCISION) & MULTS_2_9(8)(PERCISION downto 1))+signed(MULTS_2_10(8)(PERCISION) & MULTS_2_10(8)(PERCISION downto 1));
			MULTS_3_5(9)<=signed(MULTS_2_9(9)(PERCISION) & MULTS_2_9(9)(PERCISION downto 1))+signed(MULTS_2_10(9)(PERCISION) & MULTS_2_10(9)(PERCISION downto 1));
			MULTS_3_5(10)<=signed(MULTS_2_9(10)(PERCISION) & MULTS_2_9(10)(PERCISION downto 1))+signed(MULTS_2_10(10)(PERCISION) & MULTS_2_10(10)(PERCISION downto 1));
			MULTS_3_5(11)<=signed(MULTS_2_9(11)(PERCISION) & MULTS_2_9(11)(PERCISION downto 1))+signed(MULTS_2_10(11)(PERCISION) & MULTS_2_10(11)(PERCISION downto 1));
			MULTS_3_5(12)<=signed(MULTS_2_9(12)(PERCISION) & MULTS_2_9(12)(PERCISION downto 1))+signed(MULTS_2_10(12)(PERCISION) & MULTS_2_10(12)(PERCISION downto 1));
			MULTS_3_5(13)<=signed(MULTS_2_9(13)(PERCISION) & MULTS_2_9(13)(PERCISION downto 1))+signed(MULTS_2_10(13)(PERCISION) & MULTS_2_10(13)(PERCISION downto 1));
			MULTS_3_5(14)<=signed(MULTS_2_9(14)(PERCISION) & MULTS_2_9(14)(PERCISION downto 1))+signed(MULTS_2_10(14)(PERCISION) & MULTS_2_10(14)(PERCISION downto 1));
			MULTS_3_5(15)<=signed(MULTS_2_9(15)(PERCISION) & MULTS_2_9(15)(PERCISION downto 1))+signed(MULTS_2_10(15)(PERCISION) & MULTS_2_10(15)(PERCISION downto 1));
			MULTS_3_5(16)<=signed(MULTS_2_9(16)(PERCISION) & MULTS_2_9(16)(PERCISION downto 1))+signed(MULTS_2_10(16)(PERCISION) & MULTS_2_10(16)(PERCISION downto 1));
			MULTS_3_5(17)<=signed(MULTS_2_9(17)(PERCISION) & MULTS_2_9(17)(PERCISION downto 1))+signed(MULTS_2_10(17)(PERCISION) & MULTS_2_10(17)(PERCISION downto 1));
			MULTS_3_5(18)<=signed(MULTS_2_9(18)(PERCISION) & MULTS_2_9(18)(PERCISION downto 1))+signed(MULTS_2_10(18)(PERCISION) & MULTS_2_10(18)(PERCISION downto 1));
			MULTS_3_5(19)<=signed(MULTS_2_9(19)(PERCISION) & MULTS_2_9(19)(PERCISION downto 1))+signed(MULTS_2_10(19)(PERCISION) & MULTS_2_10(19)(PERCISION downto 1));
			MULTS_3_5(20)<=signed(MULTS_2_9(20)(PERCISION) & MULTS_2_9(20)(PERCISION downto 1))+signed(MULTS_2_10(20)(PERCISION) & MULTS_2_10(20)(PERCISION downto 1));
			MULTS_3_5(21)<=signed(MULTS_2_9(21)(PERCISION) & MULTS_2_9(21)(PERCISION downto 1))+signed(MULTS_2_10(21)(PERCISION) & MULTS_2_10(21)(PERCISION downto 1));
			MULTS_3_5(22)<=signed(MULTS_2_9(22)(PERCISION) & MULTS_2_9(22)(PERCISION downto 1))+signed(MULTS_2_10(22)(PERCISION) & MULTS_2_10(22)(PERCISION downto 1));
			MULTS_3_5(23)<=signed(MULTS_2_9(23)(PERCISION) & MULTS_2_9(23)(PERCISION downto 1))+signed(MULTS_2_10(23)(PERCISION) & MULTS_2_10(23)(PERCISION downto 1));
			MULTS_3_5(24)<=signed(MULTS_2_9(24)(PERCISION) & MULTS_2_9(24)(PERCISION downto 1))+signed(MULTS_2_10(24)(PERCISION) & MULTS_2_10(24)(PERCISION downto 1));
			MULTS_3_5(25)<=signed(MULTS_2_9(25)(PERCISION) & MULTS_2_9(25)(PERCISION downto 1))+signed(MULTS_2_10(25)(PERCISION) & MULTS_2_10(25)(PERCISION downto 1));
			MULTS_3_5(26)<=signed(MULTS_2_9(26)(PERCISION) & MULTS_2_9(26)(PERCISION downto 1))+signed(MULTS_2_10(26)(PERCISION) & MULTS_2_10(26)(PERCISION downto 1));
			MULTS_3_5(27)<=signed(MULTS_2_9(27)(PERCISION) & MULTS_2_9(27)(PERCISION downto 1))+signed(MULTS_2_10(27)(PERCISION) & MULTS_2_10(27)(PERCISION downto 1));
			MULTS_3_5(28)<=signed(MULTS_2_9(28)(PERCISION) & MULTS_2_9(28)(PERCISION downto 1))+signed(MULTS_2_10(28)(PERCISION) & MULTS_2_10(28)(PERCISION downto 1));
			MULTS_3_5(29)<=signed(MULTS_2_9(29)(PERCISION) & MULTS_2_9(29)(PERCISION downto 1))+signed(MULTS_2_10(29)(PERCISION) & MULTS_2_10(29)(PERCISION downto 1));
			MULTS_3_5(30)<=signed(MULTS_2_9(30)(PERCISION) & MULTS_2_9(30)(PERCISION downto 1))+signed(MULTS_2_10(30)(PERCISION) & MULTS_2_10(30)(PERCISION downto 1));
			MULTS_3_5(31)<=signed(MULTS_2_9(31)(PERCISION) & MULTS_2_9(31)(PERCISION downto 1))+signed(MULTS_2_10(31)(PERCISION) & MULTS_2_10(31)(PERCISION downto 1));
			MULTS_3_5(32)<=signed(MULTS_2_9(32)(PERCISION) & MULTS_2_9(32)(PERCISION downto 1))+signed(MULTS_2_10(32)(PERCISION) & MULTS_2_10(32)(PERCISION downto 1));
			MULTS_3_5(33)<=signed(MULTS_2_9(33)(PERCISION) & MULTS_2_9(33)(PERCISION downto 1))+signed(MULTS_2_10(33)(PERCISION) & MULTS_2_10(33)(PERCISION downto 1));
			MULTS_3_5(34)<=signed(MULTS_2_9(34)(PERCISION) & MULTS_2_9(34)(PERCISION downto 1))+signed(MULTS_2_10(34)(PERCISION) & MULTS_2_10(34)(PERCISION downto 1));
			MULTS_3_5(35)<=signed(MULTS_2_9(35)(PERCISION) & MULTS_2_9(35)(PERCISION downto 1))+signed(MULTS_2_10(35)(PERCISION) & MULTS_2_10(35)(PERCISION downto 1));
			MULTS_3_5(36)<=signed(MULTS_2_9(36)(PERCISION) & MULTS_2_9(36)(PERCISION downto 1))+signed(MULTS_2_10(36)(PERCISION) & MULTS_2_10(36)(PERCISION downto 1));
			MULTS_3_5(37)<=signed(MULTS_2_9(37)(PERCISION) & MULTS_2_9(37)(PERCISION downto 1))+signed(MULTS_2_10(37)(PERCISION) & MULTS_2_10(37)(PERCISION downto 1));
			MULTS_3_5(38)<=signed(MULTS_2_9(38)(PERCISION) & MULTS_2_9(38)(PERCISION downto 1))+signed(MULTS_2_10(38)(PERCISION) & MULTS_2_10(38)(PERCISION downto 1));
			MULTS_3_5(39)<=signed(MULTS_2_9(39)(PERCISION) & MULTS_2_9(39)(PERCISION downto 1))+signed(MULTS_2_10(39)(PERCISION) & MULTS_2_10(39)(PERCISION downto 1));
			MULTS_3_5(40)<=signed(MULTS_2_9(40)(PERCISION) & MULTS_2_9(40)(PERCISION downto 1))+signed(MULTS_2_10(40)(PERCISION) & MULTS_2_10(40)(PERCISION downto 1));
			MULTS_3_5(41)<=signed(MULTS_2_9(41)(PERCISION) & MULTS_2_9(41)(PERCISION downto 1))+signed(MULTS_2_10(41)(PERCISION) & MULTS_2_10(41)(PERCISION downto 1));
			MULTS_3_5(42)<=signed(MULTS_2_9(42)(PERCISION) & MULTS_2_9(42)(PERCISION downto 1))+signed(MULTS_2_10(42)(PERCISION) & MULTS_2_10(42)(PERCISION downto 1));
			MULTS_3_5(43)<=signed(MULTS_2_9(43)(PERCISION) & MULTS_2_9(43)(PERCISION downto 1))+signed(MULTS_2_10(43)(PERCISION) & MULTS_2_10(43)(PERCISION downto 1));
			MULTS_3_5(44)<=signed(MULTS_2_9(44)(PERCISION) & MULTS_2_9(44)(PERCISION downto 1))+signed(MULTS_2_10(44)(PERCISION) & MULTS_2_10(44)(PERCISION downto 1));
			MULTS_3_5(45)<=signed(MULTS_2_9(45)(PERCISION) & MULTS_2_9(45)(PERCISION downto 1))+signed(MULTS_2_10(45)(PERCISION) & MULTS_2_10(45)(PERCISION downto 1));
			MULTS_3_5(46)<=signed(MULTS_2_9(46)(PERCISION) & MULTS_2_9(46)(PERCISION downto 1))+signed(MULTS_2_10(46)(PERCISION) & MULTS_2_10(46)(PERCISION downto 1));
			MULTS_3_5(47)<=signed(MULTS_2_9(47)(PERCISION) & MULTS_2_9(47)(PERCISION downto 1))+signed(MULTS_2_10(47)(PERCISION) & MULTS_2_10(47)(PERCISION downto 1));
			MULTS_3_5(48)<=signed(MULTS_2_9(48)(PERCISION) & MULTS_2_9(48)(PERCISION downto 1))+signed(MULTS_2_10(48)(PERCISION) & MULTS_2_10(48)(PERCISION downto 1));
			MULTS_3_5(49)<=signed(MULTS_2_9(49)(PERCISION) & MULTS_2_9(49)(PERCISION downto 1))+signed(MULTS_2_10(49)(PERCISION) & MULTS_2_10(49)(PERCISION downto 1));
			MULTS_3_5(50)<=signed(MULTS_2_9(50)(PERCISION) & MULTS_2_9(50)(PERCISION downto 1))+signed(MULTS_2_10(50)(PERCISION) & MULTS_2_10(50)(PERCISION downto 1));
			MULTS_3_5(51)<=signed(MULTS_2_9(51)(PERCISION) & MULTS_2_9(51)(PERCISION downto 1))+signed(MULTS_2_10(51)(PERCISION) & MULTS_2_10(51)(PERCISION downto 1));
			MULTS_3_5(52)<=signed(MULTS_2_9(52)(PERCISION) & MULTS_2_9(52)(PERCISION downto 1))+signed(MULTS_2_10(52)(PERCISION) & MULTS_2_10(52)(PERCISION downto 1));
			MULTS_3_5(53)<=signed(MULTS_2_9(53)(PERCISION) & MULTS_2_9(53)(PERCISION downto 1))+signed(MULTS_2_10(53)(PERCISION) & MULTS_2_10(53)(PERCISION downto 1));
			MULTS_3_5(54)<=signed(MULTS_2_9(54)(PERCISION) & MULTS_2_9(54)(PERCISION downto 1))+signed(MULTS_2_10(54)(PERCISION) & MULTS_2_10(54)(PERCISION downto 1));
			MULTS_3_5(55)<=signed(MULTS_2_9(55)(PERCISION) & MULTS_2_9(55)(PERCISION downto 1))+signed(MULTS_2_10(55)(PERCISION) & MULTS_2_10(55)(PERCISION downto 1));
			MULTS_3_5(56)<=signed(MULTS_2_9(56)(PERCISION) & MULTS_2_9(56)(PERCISION downto 1))+signed(MULTS_2_10(56)(PERCISION) & MULTS_2_10(56)(PERCISION downto 1));
			MULTS_3_5(57)<=signed(MULTS_2_9(57)(PERCISION) & MULTS_2_9(57)(PERCISION downto 1))+signed(MULTS_2_10(57)(PERCISION) & MULTS_2_10(57)(PERCISION downto 1));
			MULTS_3_5(58)<=signed(MULTS_2_9(58)(PERCISION) & MULTS_2_9(58)(PERCISION downto 1))+signed(MULTS_2_10(58)(PERCISION) & MULTS_2_10(58)(PERCISION downto 1));
			MULTS_3_5(59)<=signed(MULTS_2_9(59)(PERCISION) & MULTS_2_9(59)(PERCISION downto 1))+signed(MULTS_2_10(59)(PERCISION) & MULTS_2_10(59)(PERCISION downto 1));
			MULTS_3_5(60)<=signed(MULTS_2_9(60)(PERCISION) & MULTS_2_9(60)(PERCISION downto 1))+signed(MULTS_2_10(60)(PERCISION) & MULTS_2_10(60)(PERCISION downto 1));
			MULTS_3_5(61)<=signed(MULTS_2_9(61)(PERCISION) & MULTS_2_9(61)(PERCISION downto 1))+signed(MULTS_2_10(61)(PERCISION) & MULTS_2_10(61)(PERCISION downto 1));
			MULTS_3_5(62)<=signed(MULTS_2_9(62)(PERCISION) & MULTS_2_9(62)(PERCISION downto 1))+signed(MULTS_2_10(62)(PERCISION) & MULTS_2_10(62)(PERCISION downto 1));
			MULTS_3_5(63)<=signed(MULTS_2_9(63)(PERCISION) & MULTS_2_9(63)(PERCISION downto 1))+signed(MULTS_2_10(63)(PERCISION) & MULTS_2_10(63)(PERCISION downto 1));
			MULTS_3_5(64)<=signed(MULTS_2_9(64)(PERCISION) & MULTS_2_9(64)(PERCISION downto 1))+signed(MULTS_2_10(64)(PERCISION) & MULTS_2_10(64)(PERCISION downto 1));
			MULTS_3_5(65)<=signed(MULTS_2_9(65)(PERCISION) & MULTS_2_9(65)(PERCISION downto 1))+signed(MULTS_2_10(65)(PERCISION) & MULTS_2_10(65)(PERCISION downto 1));
			MULTS_3_5(66)<=signed(MULTS_2_9(66)(PERCISION) & MULTS_2_9(66)(PERCISION downto 1))+signed(MULTS_2_10(66)(PERCISION) & MULTS_2_10(66)(PERCISION downto 1));
			MULTS_3_5(67)<=signed(MULTS_2_9(67)(PERCISION) & MULTS_2_9(67)(PERCISION downto 1))+signed(MULTS_2_10(67)(PERCISION) & MULTS_2_10(67)(PERCISION downto 1));
			MULTS_3_5(68)<=signed(MULTS_2_9(68)(PERCISION) & MULTS_2_9(68)(PERCISION downto 1))+signed(MULTS_2_10(68)(PERCISION) & MULTS_2_10(68)(PERCISION downto 1));
			MULTS_3_5(69)<=signed(MULTS_2_9(69)(PERCISION) & MULTS_2_9(69)(PERCISION downto 1))+signed(MULTS_2_10(69)(PERCISION) & MULTS_2_10(69)(PERCISION downto 1));
			MULTS_3_5(70)<=signed(MULTS_2_9(70)(PERCISION) & MULTS_2_9(70)(PERCISION downto 1))+signed(MULTS_2_10(70)(PERCISION) & MULTS_2_10(70)(PERCISION downto 1));
			MULTS_3_5(71)<=signed(MULTS_2_9(71)(PERCISION) & MULTS_2_9(71)(PERCISION downto 1))+signed(MULTS_2_10(71)(PERCISION) & MULTS_2_10(71)(PERCISION downto 1));
			MULTS_3_5(72)<=signed(MULTS_2_9(72)(PERCISION) & MULTS_2_9(72)(PERCISION downto 1))+signed(MULTS_2_10(72)(PERCISION) & MULTS_2_10(72)(PERCISION downto 1));
			MULTS_3_5(73)<=signed(MULTS_2_9(73)(PERCISION) & MULTS_2_9(73)(PERCISION downto 1))+signed(MULTS_2_10(73)(PERCISION) & MULTS_2_10(73)(PERCISION downto 1));
			MULTS_3_5(74)<=signed(MULTS_2_9(74)(PERCISION) & MULTS_2_9(74)(PERCISION downto 1))+signed(MULTS_2_10(74)(PERCISION) & MULTS_2_10(74)(PERCISION downto 1));
			MULTS_3_5(75)<=signed(MULTS_2_9(75)(PERCISION) & MULTS_2_9(75)(PERCISION downto 1))+signed(MULTS_2_10(75)(PERCISION) & MULTS_2_10(75)(PERCISION downto 1));
			MULTS_3_5(76)<=signed(MULTS_2_9(76)(PERCISION) & MULTS_2_9(76)(PERCISION downto 1))+signed(MULTS_2_10(76)(PERCISION) & MULTS_2_10(76)(PERCISION downto 1));
			MULTS_3_5(77)<=signed(MULTS_2_9(77)(PERCISION) & MULTS_2_9(77)(PERCISION downto 1))+signed(MULTS_2_10(77)(PERCISION) & MULTS_2_10(77)(PERCISION downto 1));
			MULTS_3_5(78)<=signed(MULTS_2_9(78)(PERCISION) & MULTS_2_9(78)(PERCISION downto 1))+signed(MULTS_2_10(78)(PERCISION) & MULTS_2_10(78)(PERCISION downto 1));
			MULTS_3_5(79)<=signed(MULTS_2_9(79)(PERCISION) & MULTS_2_9(79)(PERCISION downto 1))+signed(MULTS_2_10(79)(PERCISION) & MULTS_2_10(79)(PERCISION downto 1));
			MULTS_3_5(80)<=signed(MULTS_2_9(80)(PERCISION) & MULTS_2_9(80)(PERCISION downto 1))+signed(MULTS_2_10(80)(PERCISION) & MULTS_2_10(80)(PERCISION downto 1));
			MULTS_3_5(81)<=signed(MULTS_2_9(81)(PERCISION) & MULTS_2_9(81)(PERCISION downto 1))+signed(MULTS_2_10(81)(PERCISION) & MULTS_2_10(81)(PERCISION downto 1));
			MULTS_3_5(82)<=signed(MULTS_2_9(82)(PERCISION) & MULTS_2_9(82)(PERCISION downto 1))+signed(MULTS_2_10(82)(PERCISION) & MULTS_2_10(82)(PERCISION downto 1));
			MULTS_3_5(83)<=signed(MULTS_2_9(83)(PERCISION) & MULTS_2_9(83)(PERCISION downto 1))+signed(MULTS_2_10(83)(PERCISION) & MULTS_2_10(83)(PERCISION downto 1));

			MULTS_3_6(0)<=signed(MULTS_2_11(0)(PERCISION) & MULTS_2_11(0)(PERCISION downto 1))+signed(MULTS_2_12(0)(PERCISION) & MULTS_2_12(0)(PERCISION downto 1));
			MULTS_3_6(1)<=signed(MULTS_2_11(1)(PERCISION) & MULTS_2_11(1)(PERCISION downto 1))+signed(MULTS_2_12(1)(PERCISION) & MULTS_2_12(1)(PERCISION downto 1));
			MULTS_3_6(2)<=signed(MULTS_2_11(2)(PERCISION) & MULTS_2_11(2)(PERCISION downto 1))+signed(MULTS_2_12(2)(PERCISION) & MULTS_2_12(2)(PERCISION downto 1));
			MULTS_3_6(3)<=signed(MULTS_2_11(3)(PERCISION) & MULTS_2_11(3)(PERCISION downto 1))+signed(MULTS_2_12(3)(PERCISION) & MULTS_2_12(3)(PERCISION downto 1));
			MULTS_3_6(4)<=signed(MULTS_2_11(4)(PERCISION) & MULTS_2_11(4)(PERCISION downto 1))+signed(MULTS_2_12(4)(PERCISION) & MULTS_2_12(4)(PERCISION downto 1));
			MULTS_3_6(5)<=signed(MULTS_2_11(5)(PERCISION) & MULTS_2_11(5)(PERCISION downto 1))+signed(MULTS_2_12(5)(PERCISION) & MULTS_2_12(5)(PERCISION downto 1));
			MULTS_3_6(6)<=signed(MULTS_2_11(6)(PERCISION) & MULTS_2_11(6)(PERCISION downto 1))+signed(MULTS_2_12(6)(PERCISION) & MULTS_2_12(6)(PERCISION downto 1));
			MULTS_3_6(7)<=signed(MULTS_2_11(7)(PERCISION) & MULTS_2_11(7)(PERCISION downto 1))+signed(MULTS_2_12(7)(PERCISION) & MULTS_2_12(7)(PERCISION downto 1));
			MULTS_3_6(8)<=signed(MULTS_2_11(8)(PERCISION) & MULTS_2_11(8)(PERCISION downto 1))+signed(MULTS_2_12(8)(PERCISION) & MULTS_2_12(8)(PERCISION downto 1));
			MULTS_3_6(9)<=signed(MULTS_2_11(9)(PERCISION) & MULTS_2_11(9)(PERCISION downto 1))+signed(MULTS_2_12(9)(PERCISION) & MULTS_2_12(9)(PERCISION downto 1));
			MULTS_3_6(10)<=signed(MULTS_2_11(10)(PERCISION) & MULTS_2_11(10)(PERCISION downto 1))+signed(MULTS_2_12(10)(PERCISION) & MULTS_2_12(10)(PERCISION downto 1));
			MULTS_3_6(11)<=signed(MULTS_2_11(11)(PERCISION) & MULTS_2_11(11)(PERCISION downto 1))+signed(MULTS_2_12(11)(PERCISION) & MULTS_2_12(11)(PERCISION downto 1));
			MULTS_3_6(12)<=signed(MULTS_2_11(12)(PERCISION) & MULTS_2_11(12)(PERCISION downto 1))+signed(MULTS_2_12(12)(PERCISION) & MULTS_2_12(12)(PERCISION downto 1));
			MULTS_3_6(13)<=signed(MULTS_2_11(13)(PERCISION) & MULTS_2_11(13)(PERCISION downto 1))+signed(MULTS_2_12(13)(PERCISION) & MULTS_2_12(13)(PERCISION downto 1));
			MULTS_3_6(14)<=signed(MULTS_2_11(14)(PERCISION) & MULTS_2_11(14)(PERCISION downto 1))+signed(MULTS_2_12(14)(PERCISION) & MULTS_2_12(14)(PERCISION downto 1));
			MULTS_3_6(15)<=signed(MULTS_2_11(15)(PERCISION) & MULTS_2_11(15)(PERCISION downto 1))+signed(MULTS_2_12(15)(PERCISION) & MULTS_2_12(15)(PERCISION downto 1));
			MULTS_3_6(16)<=signed(MULTS_2_11(16)(PERCISION) & MULTS_2_11(16)(PERCISION downto 1))+signed(MULTS_2_12(16)(PERCISION) & MULTS_2_12(16)(PERCISION downto 1));
			MULTS_3_6(17)<=signed(MULTS_2_11(17)(PERCISION) & MULTS_2_11(17)(PERCISION downto 1))+signed(MULTS_2_12(17)(PERCISION) & MULTS_2_12(17)(PERCISION downto 1));
			MULTS_3_6(18)<=signed(MULTS_2_11(18)(PERCISION) & MULTS_2_11(18)(PERCISION downto 1))+signed(MULTS_2_12(18)(PERCISION) & MULTS_2_12(18)(PERCISION downto 1));
			MULTS_3_6(19)<=signed(MULTS_2_11(19)(PERCISION) & MULTS_2_11(19)(PERCISION downto 1))+signed(MULTS_2_12(19)(PERCISION) & MULTS_2_12(19)(PERCISION downto 1));
			MULTS_3_6(20)<=signed(MULTS_2_11(20)(PERCISION) & MULTS_2_11(20)(PERCISION downto 1))+signed(MULTS_2_12(20)(PERCISION) & MULTS_2_12(20)(PERCISION downto 1));
			MULTS_3_6(21)<=signed(MULTS_2_11(21)(PERCISION) & MULTS_2_11(21)(PERCISION downto 1))+signed(MULTS_2_12(21)(PERCISION) & MULTS_2_12(21)(PERCISION downto 1));
			MULTS_3_6(22)<=signed(MULTS_2_11(22)(PERCISION) & MULTS_2_11(22)(PERCISION downto 1))+signed(MULTS_2_12(22)(PERCISION) & MULTS_2_12(22)(PERCISION downto 1));
			MULTS_3_6(23)<=signed(MULTS_2_11(23)(PERCISION) & MULTS_2_11(23)(PERCISION downto 1))+signed(MULTS_2_12(23)(PERCISION) & MULTS_2_12(23)(PERCISION downto 1));
			MULTS_3_6(24)<=signed(MULTS_2_11(24)(PERCISION) & MULTS_2_11(24)(PERCISION downto 1))+signed(MULTS_2_12(24)(PERCISION) & MULTS_2_12(24)(PERCISION downto 1));
			MULTS_3_6(25)<=signed(MULTS_2_11(25)(PERCISION) & MULTS_2_11(25)(PERCISION downto 1))+signed(MULTS_2_12(25)(PERCISION) & MULTS_2_12(25)(PERCISION downto 1));
			MULTS_3_6(26)<=signed(MULTS_2_11(26)(PERCISION) & MULTS_2_11(26)(PERCISION downto 1))+signed(MULTS_2_12(26)(PERCISION) & MULTS_2_12(26)(PERCISION downto 1));
			MULTS_3_6(27)<=signed(MULTS_2_11(27)(PERCISION) & MULTS_2_11(27)(PERCISION downto 1))+signed(MULTS_2_12(27)(PERCISION) & MULTS_2_12(27)(PERCISION downto 1));
			MULTS_3_6(28)<=signed(MULTS_2_11(28)(PERCISION) & MULTS_2_11(28)(PERCISION downto 1))+signed(MULTS_2_12(28)(PERCISION) & MULTS_2_12(28)(PERCISION downto 1));
			MULTS_3_6(29)<=signed(MULTS_2_11(29)(PERCISION) & MULTS_2_11(29)(PERCISION downto 1))+signed(MULTS_2_12(29)(PERCISION) & MULTS_2_12(29)(PERCISION downto 1));
			MULTS_3_6(30)<=signed(MULTS_2_11(30)(PERCISION) & MULTS_2_11(30)(PERCISION downto 1))+signed(MULTS_2_12(30)(PERCISION) & MULTS_2_12(30)(PERCISION downto 1));
			MULTS_3_6(31)<=signed(MULTS_2_11(31)(PERCISION) & MULTS_2_11(31)(PERCISION downto 1))+signed(MULTS_2_12(31)(PERCISION) & MULTS_2_12(31)(PERCISION downto 1));
			MULTS_3_6(32)<=signed(MULTS_2_11(32)(PERCISION) & MULTS_2_11(32)(PERCISION downto 1))+signed(MULTS_2_12(32)(PERCISION) & MULTS_2_12(32)(PERCISION downto 1));
			MULTS_3_6(33)<=signed(MULTS_2_11(33)(PERCISION) & MULTS_2_11(33)(PERCISION downto 1))+signed(MULTS_2_12(33)(PERCISION) & MULTS_2_12(33)(PERCISION downto 1));
			MULTS_3_6(34)<=signed(MULTS_2_11(34)(PERCISION) & MULTS_2_11(34)(PERCISION downto 1))+signed(MULTS_2_12(34)(PERCISION) & MULTS_2_12(34)(PERCISION downto 1));
			MULTS_3_6(35)<=signed(MULTS_2_11(35)(PERCISION) & MULTS_2_11(35)(PERCISION downto 1))+signed(MULTS_2_12(35)(PERCISION) & MULTS_2_12(35)(PERCISION downto 1));
			MULTS_3_6(36)<=signed(MULTS_2_11(36)(PERCISION) & MULTS_2_11(36)(PERCISION downto 1))+signed(MULTS_2_12(36)(PERCISION) & MULTS_2_12(36)(PERCISION downto 1));
			MULTS_3_6(37)<=signed(MULTS_2_11(37)(PERCISION) & MULTS_2_11(37)(PERCISION downto 1))+signed(MULTS_2_12(37)(PERCISION) & MULTS_2_12(37)(PERCISION downto 1));
			MULTS_3_6(38)<=signed(MULTS_2_11(38)(PERCISION) & MULTS_2_11(38)(PERCISION downto 1))+signed(MULTS_2_12(38)(PERCISION) & MULTS_2_12(38)(PERCISION downto 1));
			MULTS_3_6(39)<=signed(MULTS_2_11(39)(PERCISION) & MULTS_2_11(39)(PERCISION downto 1))+signed(MULTS_2_12(39)(PERCISION) & MULTS_2_12(39)(PERCISION downto 1));
			MULTS_3_6(40)<=signed(MULTS_2_11(40)(PERCISION) & MULTS_2_11(40)(PERCISION downto 1))+signed(MULTS_2_12(40)(PERCISION) & MULTS_2_12(40)(PERCISION downto 1));
			MULTS_3_6(41)<=signed(MULTS_2_11(41)(PERCISION) & MULTS_2_11(41)(PERCISION downto 1))+signed(MULTS_2_12(41)(PERCISION) & MULTS_2_12(41)(PERCISION downto 1));
			MULTS_3_6(42)<=signed(MULTS_2_11(42)(PERCISION) & MULTS_2_11(42)(PERCISION downto 1))+signed(MULTS_2_12(42)(PERCISION) & MULTS_2_12(42)(PERCISION downto 1));
			MULTS_3_6(43)<=signed(MULTS_2_11(43)(PERCISION) & MULTS_2_11(43)(PERCISION downto 1))+signed(MULTS_2_12(43)(PERCISION) & MULTS_2_12(43)(PERCISION downto 1));
			MULTS_3_6(44)<=signed(MULTS_2_11(44)(PERCISION) & MULTS_2_11(44)(PERCISION downto 1))+signed(MULTS_2_12(44)(PERCISION) & MULTS_2_12(44)(PERCISION downto 1));
			MULTS_3_6(45)<=signed(MULTS_2_11(45)(PERCISION) & MULTS_2_11(45)(PERCISION downto 1))+signed(MULTS_2_12(45)(PERCISION) & MULTS_2_12(45)(PERCISION downto 1));
			MULTS_3_6(46)<=signed(MULTS_2_11(46)(PERCISION) & MULTS_2_11(46)(PERCISION downto 1))+signed(MULTS_2_12(46)(PERCISION) & MULTS_2_12(46)(PERCISION downto 1));
			MULTS_3_6(47)<=signed(MULTS_2_11(47)(PERCISION) & MULTS_2_11(47)(PERCISION downto 1))+signed(MULTS_2_12(47)(PERCISION) & MULTS_2_12(47)(PERCISION downto 1));
			MULTS_3_6(48)<=signed(MULTS_2_11(48)(PERCISION) & MULTS_2_11(48)(PERCISION downto 1))+signed(MULTS_2_12(48)(PERCISION) & MULTS_2_12(48)(PERCISION downto 1));
			MULTS_3_6(49)<=signed(MULTS_2_11(49)(PERCISION) & MULTS_2_11(49)(PERCISION downto 1))+signed(MULTS_2_12(49)(PERCISION) & MULTS_2_12(49)(PERCISION downto 1));
			MULTS_3_6(50)<=signed(MULTS_2_11(50)(PERCISION) & MULTS_2_11(50)(PERCISION downto 1))+signed(MULTS_2_12(50)(PERCISION) & MULTS_2_12(50)(PERCISION downto 1));
			MULTS_3_6(51)<=signed(MULTS_2_11(51)(PERCISION) & MULTS_2_11(51)(PERCISION downto 1))+signed(MULTS_2_12(51)(PERCISION) & MULTS_2_12(51)(PERCISION downto 1));
			MULTS_3_6(52)<=signed(MULTS_2_11(52)(PERCISION) & MULTS_2_11(52)(PERCISION downto 1))+signed(MULTS_2_12(52)(PERCISION) & MULTS_2_12(52)(PERCISION downto 1));
			MULTS_3_6(53)<=signed(MULTS_2_11(53)(PERCISION) & MULTS_2_11(53)(PERCISION downto 1))+signed(MULTS_2_12(53)(PERCISION) & MULTS_2_12(53)(PERCISION downto 1));
			MULTS_3_6(54)<=signed(MULTS_2_11(54)(PERCISION) & MULTS_2_11(54)(PERCISION downto 1))+signed(MULTS_2_12(54)(PERCISION) & MULTS_2_12(54)(PERCISION downto 1));
			MULTS_3_6(55)<=signed(MULTS_2_11(55)(PERCISION) & MULTS_2_11(55)(PERCISION downto 1))+signed(MULTS_2_12(55)(PERCISION) & MULTS_2_12(55)(PERCISION downto 1));
			MULTS_3_6(56)<=signed(MULTS_2_11(56)(PERCISION) & MULTS_2_11(56)(PERCISION downto 1))+signed(MULTS_2_12(56)(PERCISION) & MULTS_2_12(56)(PERCISION downto 1));
			MULTS_3_6(57)<=signed(MULTS_2_11(57)(PERCISION) & MULTS_2_11(57)(PERCISION downto 1))+signed(MULTS_2_12(57)(PERCISION) & MULTS_2_12(57)(PERCISION downto 1));
			MULTS_3_6(58)<=signed(MULTS_2_11(58)(PERCISION) & MULTS_2_11(58)(PERCISION downto 1))+signed(MULTS_2_12(58)(PERCISION) & MULTS_2_12(58)(PERCISION downto 1));
			MULTS_3_6(59)<=signed(MULTS_2_11(59)(PERCISION) & MULTS_2_11(59)(PERCISION downto 1))+signed(MULTS_2_12(59)(PERCISION) & MULTS_2_12(59)(PERCISION downto 1));
			MULTS_3_6(60)<=signed(MULTS_2_11(60)(PERCISION) & MULTS_2_11(60)(PERCISION downto 1))+signed(MULTS_2_12(60)(PERCISION) & MULTS_2_12(60)(PERCISION downto 1));
			MULTS_3_6(61)<=signed(MULTS_2_11(61)(PERCISION) & MULTS_2_11(61)(PERCISION downto 1))+signed(MULTS_2_12(61)(PERCISION) & MULTS_2_12(61)(PERCISION downto 1));
			MULTS_3_6(62)<=signed(MULTS_2_11(62)(PERCISION) & MULTS_2_11(62)(PERCISION downto 1))+signed(MULTS_2_12(62)(PERCISION) & MULTS_2_12(62)(PERCISION downto 1));
			MULTS_3_6(63)<=signed(MULTS_2_11(63)(PERCISION) & MULTS_2_11(63)(PERCISION downto 1))+signed(MULTS_2_12(63)(PERCISION) & MULTS_2_12(63)(PERCISION downto 1));
			MULTS_3_6(64)<=signed(MULTS_2_11(64)(PERCISION) & MULTS_2_11(64)(PERCISION downto 1))+signed(MULTS_2_12(64)(PERCISION) & MULTS_2_12(64)(PERCISION downto 1));
			MULTS_3_6(65)<=signed(MULTS_2_11(65)(PERCISION) & MULTS_2_11(65)(PERCISION downto 1))+signed(MULTS_2_12(65)(PERCISION) & MULTS_2_12(65)(PERCISION downto 1));
			MULTS_3_6(66)<=signed(MULTS_2_11(66)(PERCISION) & MULTS_2_11(66)(PERCISION downto 1))+signed(MULTS_2_12(66)(PERCISION) & MULTS_2_12(66)(PERCISION downto 1));
			MULTS_3_6(67)<=signed(MULTS_2_11(67)(PERCISION) & MULTS_2_11(67)(PERCISION downto 1))+signed(MULTS_2_12(67)(PERCISION) & MULTS_2_12(67)(PERCISION downto 1));
			MULTS_3_6(68)<=signed(MULTS_2_11(68)(PERCISION) & MULTS_2_11(68)(PERCISION downto 1))+signed(MULTS_2_12(68)(PERCISION) & MULTS_2_12(68)(PERCISION downto 1));
			MULTS_3_6(69)<=signed(MULTS_2_11(69)(PERCISION) & MULTS_2_11(69)(PERCISION downto 1))+signed(MULTS_2_12(69)(PERCISION) & MULTS_2_12(69)(PERCISION downto 1));
			MULTS_3_6(70)<=signed(MULTS_2_11(70)(PERCISION) & MULTS_2_11(70)(PERCISION downto 1))+signed(MULTS_2_12(70)(PERCISION) & MULTS_2_12(70)(PERCISION downto 1));
			MULTS_3_6(71)<=signed(MULTS_2_11(71)(PERCISION) & MULTS_2_11(71)(PERCISION downto 1))+signed(MULTS_2_12(71)(PERCISION) & MULTS_2_12(71)(PERCISION downto 1));
			MULTS_3_6(72)<=signed(MULTS_2_11(72)(PERCISION) & MULTS_2_11(72)(PERCISION downto 1))+signed(MULTS_2_12(72)(PERCISION) & MULTS_2_12(72)(PERCISION downto 1));
			MULTS_3_6(73)<=signed(MULTS_2_11(73)(PERCISION) & MULTS_2_11(73)(PERCISION downto 1))+signed(MULTS_2_12(73)(PERCISION) & MULTS_2_12(73)(PERCISION downto 1));
			MULTS_3_6(74)<=signed(MULTS_2_11(74)(PERCISION) & MULTS_2_11(74)(PERCISION downto 1))+signed(MULTS_2_12(74)(PERCISION) & MULTS_2_12(74)(PERCISION downto 1));
			MULTS_3_6(75)<=signed(MULTS_2_11(75)(PERCISION) & MULTS_2_11(75)(PERCISION downto 1))+signed(MULTS_2_12(75)(PERCISION) & MULTS_2_12(75)(PERCISION downto 1));
			MULTS_3_6(76)<=signed(MULTS_2_11(76)(PERCISION) & MULTS_2_11(76)(PERCISION downto 1))+signed(MULTS_2_12(76)(PERCISION) & MULTS_2_12(76)(PERCISION downto 1));
			MULTS_3_6(77)<=signed(MULTS_2_11(77)(PERCISION) & MULTS_2_11(77)(PERCISION downto 1))+signed(MULTS_2_12(77)(PERCISION) & MULTS_2_12(77)(PERCISION downto 1));
			MULTS_3_6(78)<=signed(MULTS_2_11(78)(PERCISION) & MULTS_2_11(78)(PERCISION downto 1))+signed(MULTS_2_12(78)(PERCISION) & MULTS_2_12(78)(PERCISION downto 1));
			MULTS_3_6(79)<=signed(MULTS_2_11(79)(PERCISION) & MULTS_2_11(79)(PERCISION downto 1))+signed(MULTS_2_12(79)(PERCISION) & MULTS_2_12(79)(PERCISION downto 1));
			MULTS_3_6(80)<=signed(MULTS_2_11(80)(PERCISION) & MULTS_2_11(80)(PERCISION downto 1))+signed(MULTS_2_12(80)(PERCISION) & MULTS_2_12(80)(PERCISION downto 1));
			MULTS_3_6(81)<=signed(MULTS_2_11(81)(PERCISION) & MULTS_2_11(81)(PERCISION downto 1))+signed(MULTS_2_12(81)(PERCISION) & MULTS_2_12(81)(PERCISION downto 1));
			MULTS_3_6(82)<=signed(MULTS_2_11(82)(PERCISION) & MULTS_2_11(82)(PERCISION downto 1))+signed(MULTS_2_12(82)(PERCISION) & MULTS_2_12(82)(PERCISION downto 1));
			MULTS_3_6(83)<=signed(MULTS_2_11(83)(PERCISION) & MULTS_2_11(83)(PERCISION downto 1))+signed(MULTS_2_12(83)(PERCISION) & MULTS_2_12(83)(PERCISION downto 1));

			MULTS_3_7(0)<=signed(MULTS_2_13(0)(PERCISION) & MULTS_2_13(0)(PERCISION downto 1))+signed(MULTS_2_14(0)(PERCISION) & MULTS_2_14(0)(PERCISION downto 1));
			MULTS_3_7(1)<=signed(MULTS_2_13(1)(PERCISION) & MULTS_2_13(1)(PERCISION downto 1))+signed(MULTS_2_14(1)(PERCISION) & MULTS_2_14(1)(PERCISION downto 1));
			MULTS_3_7(2)<=signed(MULTS_2_13(2)(PERCISION) & MULTS_2_13(2)(PERCISION downto 1))+signed(MULTS_2_14(2)(PERCISION) & MULTS_2_14(2)(PERCISION downto 1));
			MULTS_3_7(3)<=signed(MULTS_2_13(3)(PERCISION) & MULTS_2_13(3)(PERCISION downto 1))+signed(MULTS_2_14(3)(PERCISION) & MULTS_2_14(3)(PERCISION downto 1));
			MULTS_3_7(4)<=signed(MULTS_2_13(4)(PERCISION) & MULTS_2_13(4)(PERCISION downto 1))+signed(MULTS_2_14(4)(PERCISION) & MULTS_2_14(4)(PERCISION downto 1));
			MULTS_3_7(5)<=signed(MULTS_2_13(5)(PERCISION) & MULTS_2_13(5)(PERCISION downto 1))+signed(MULTS_2_14(5)(PERCISION) & MULTS_2_14(5)(PERCISION downto 1));
			MULTS_3_7(6)<=signed(MULTS_2_13(6)(PERCISION) & MULTS_2_13(6)(PERCISION downto 1))+signed(MULTS_2_14(6)(PERCISION) & MULTS_2_14(6)(PERCISION downto 1));
			MULTS_3_7(7)<=signed(MULTS_2_13(7)(PERCISION) & MULTS_2_13(7)(PERCISION downto 1))+signed(MULTS_2_14(7)(PERCISION) & MULTS_2_14(7)(PERCISION downto 1));
			MULTS_3_7(8)<=signed(MULTS_2_13(8)(PERCISION) & MULTS_2_13(8)(PERCISION downto 1))+signed(MULTS_2_14(8)(PERCISION) & MULTS_2_14(8)(PERCISION downto 1));
			MULTS_3_7(9)<=signed(MULTS_2_13(9)(PERCISION) & MULTS_2_13(9)(PERCISION downto 1))+signed(MULTS_2_14(9)(PERCISION) & MULTS_2_14(9)(PERCISION downto 1));
			MULTS_3_7(10)<=signed(MULTS_2_13(10)(PERCISION) & MULTS_2_13(10)(PERCISION downto 1))+signed(MULTS_2_14(10)(PERCISION) & MULTS_2_14(10)(PERCISION downto 1));
			MULTS_3_7(11)<=signed(MULTS_2_13(11)(PERCISION) & MULTS_2_13(11)(PERCISION downto 1))+signed(MULTS_2_14(11)(PERCISION) & MULTS_2_14(11)(PERCISION downto 1));
			MULTS_3_7(12)<=signed(MULTS_2_13(12)(PERCISION) & MULTS_2_13(12)(PERCISION downto 1))+signed(MULTS_2_14(12)(PERCISION) & MULTS_2_14(12)(PERCISION downto 1));
			MULTS_3_7(13)<=signed(MULTS_2_13(13)(PERCISION) & MULTS_2_13(13)(PERCISION downto 1))+signed(MULTS_2_14(13)(PERCISION) & MULTS_2_14(13)(PERCISION downto 1));
			MULTS_3_7(14)<=signed(MULTS_2_13(14)(PERCISION) & MULTS_2_13(14)(PERCISION downto 1))+signed(MULTS_2_14(14)(PERCISION) & MULTS_2_14(14)(PERCISION downto 1));
			MULTS_3_7(15)<=signed(MULTS_2_13(15)(PERCISION) & MULTS_2_13(15)(PERCISION downto 1))+signed(MULTS_2_14(15)(PERCISION) & MULTS_2_14(15)(PERCISION downto 1));
			MULTS_3_7(16)<=signed(MULTS_2_13(16)(PERCISION) & MULTS_2_13(16)(PERCISION downto 1))+signed(MULTS_2_14(16)(PERCISION) & MULTS_2_14(16)(PERCISION downto 1));
			MULTS_3_7(17)<=signed(MULTS_2_13(17)(PERCISION) & MULTS_2_13(17)(PERCISION downto 1))+signed(MULTS_2_14(17)(PERCISION) & MULTS_2_14(17)(PERCISION downto 1));
			MULTS_3_7(18)<=signed(MULTS_2_13(18)(PERCISION) & MULTS_2_13(18)(PERCISION downto 1))+signed(MULTS_2_14(18)(PERCISION) & MULTS_2_14(18)(PERCISION downto 1));
			MULTS_3_7(19)<=signed(MULTS_2_13(19)(PERCISION) & MULTS_2_13(19)(PERCISION downto 1))+signed(MULTS_2_14(19)(PERCISION) & MULTS_2_14(19)(PERCISION downto 1));
			MULTS_3_7(20)<=signed(MULTS_2_13(20)(PERCISION) & MULTS_2_13(20)(PERCISION downto 1))+signed(MULTS_2_14(20)(PERCISION) & MULTS_2_14(20)(PERCISION downto 1));
			MULTS_3_7(21)<=signed(MULTS_2_13(21)(PERCISION) & MULTS_2_13(21)(PERCISION downto 1))+signed(MULTS_2_14(21)(PERCISION) & MULTS_2_14(21)(PERCISION downto 1));
			MULTS_3_7(22)<=signed(MULTS_2_13(22)(PERCISION) & MULTS_2_13(22)(PERCISION downto 1))+signed(MULTS_2_14(22)(PERCISION) & MULTS_2_14(22)(PERCISION downto 1));
			MULTS_3_7(23)<=signed(MULTS_2_13(23)(PERCISION) & MULTS_2_13(23)(PERCISION downto 1))+signed(MULTS_2_14(23)(PERCISION) & MULTS_2_14(23)(PERCISION downto 1));
			MULTS_3_7(24)<=signed(MULTS_2_13(24)(PERCISION) & MULTS_2_13(24)(PERCISION downto 1))+signed(MULTS_2_14(24)(PERCISION) & MULTS_2_14(24)(PERCISION downto 1));
			MULTS_3_7(25)<=signed(MULTS_2_13(25)(PERCISION) & MULTS_2_13(25)(PERCISION downto 1))+signed(MULTS_2_14(25)(PERCISION) & MULTS_2_14(25)(PERCISION downto 1));
			MULTS_3_7(26)<=signed(MULTS_2_13(26)(PERCISION) & MULTS_2_13(26)(PERCISION downto 1))+signed(MULTS_2_14(26)(PERCISION) & MULTS_2_14(26)(PERCISION downto 1));
			MULTS_3_7(27)<=signed(MULTS_2_13(27)(PERCISION) & MULTS_2_13(27)(PERCISION downto 1))+signed(MULTS_2_14(27)(PERCISION) & MULTS_2_14(27)(PERCISION downto 1));
			MULTS_3_7(28)<=signed(MULTS_2_13(28)(PERCISION) & MULTS_2_13(28)(PERCISION downto 1))+signed(MULTS_2_14(28)(PERCISION) & MULTS_2_14(28)(PERCISION downto 1));
			MULTS_3_7(29)<=signed(MULTS_2_13(29)(PERCISION) & MULTS_2_13(29)(PERCISION downto 1))+signed(MULTS_2_14(29)(PERCISION) & MULTS_2_14(29)(PERCISION downto 1));
			MULTS_3_7(30)<=signed(MULTS_2_13(30)(PERCISION) & MULTS_2_13(30)(PERCISION downto 1))+signed(MULTS_2_14(30)(PERCISION) & MULTS_2_14(30)(PERCISION downto 1));
			MULTS_3_7(31)<=signed(MULTS_2_13(31)(PERCISION) & MULTS_2_13(31)(PERCISION downto 1))+signed(MULTS_2_14(31)(PERCISION) & MULTS_2_14(31)(PERCISION downto 1));
			MULTS_3_7(32)<=signed(MULTS_2_13(32)(PERCISION) & MULTS_2_13(32)(PERCISION downto 1))+signed(MULTS_2_14(32)(PERCISION) & MULTS_2_14(32)(PERCISION downto 1));
			MULTS_3_7(33)<=signed(MULTS_2_13(33)(PERCISION) & MULTS_2_13(33)(PERCISION downto 1))+signed(MULTS_2_14(33)(PERCISION) & MULTS_2_14(33)(PERCISION downto 1));
			MULTS_3_7(34)<=signed(MULTS_2_13(34)(PERCISION) & MULTS_2_13(34)(PERCISION downto 1))+signed(MULTS_2_14(34)(PERCISION) & MULTS_2_14(34)(PERCISION downto 1));
			MULTS_3_7(35)<=signed(MULTS_2_13(35)(PERCISION) & MULTS_2_13(35)(PERCISION downto 1))+signed(MULTS_2_14(35)(PERCISION) & MULTS_2_14(35)(PERCISION downto 1));
			MULTS_3_7(36)<=signed(MULTS_2_13(36)(PERCISION) & MULTS_2_13(36)(PERCISION downto 1))+signed(MULTS_2_14(36)(PERCISION) & MULTS_2_14(36)(PERCISION downto 1));
			MULTS_3_7(37)<=signed(MULTS_2_13(37)(PERCISION) & MULTS_2_13(37)(PERCISION downto 1))+signed(MULTS_2_14(37)(PERCISION) & MULTS_2_14(37)(PERCISION downto 1));
			MULTS_3_7(38)<=signed(MULTS_2_13(38)(PERCISION) & MULTS_2_13(38)(PERCISION downto 1))+signed(MULTS_2_14(38)(PERCISION) & MULTS_2_14(38)(PERCISION downto 1));
			MULTS_3_7(39)<=signed(MULTS_2_13(39)(PERCISION) & MULTS_2_13(39)(PERCISION downto 1))+signed(MULTS_2_14(39)(PERCISION) & MULTS_2_14(39)(PERCISION downto 1));
			MULTS_3_7(40)<=signed(MULTS_2_13(40)(PERCISION) & MULTS_2_13(40)(PERCISION downto 1))+signed(MULTS_2_14(40)(PERCISION) & MULTS_2_14(40)(PERCISION downto 1));
			MULTS_3_7(41)<=signed(MULTS_2_13(41)(PERCISION) & MULTS_2_13(41)(PERCISION downto 1))+signed(MULTS_2_14(41)(PERCISION) & MULTS_2_14(41)(PERCISION downto 1));
			MULTS_3_7(42)<=signed(MULTS_2_13(42)(PERCISION) & MULTS_2_13(42)(PERCISION downto 1))+signed(MULTS_2_14(42)(PERCISION) & MULTS_2_14(42)(PERCISION downto 1));
			MULTS_3_7(43)<=signed(MULTS_2_13(43)(PERCISION) & MULTS_2_13(43)(PERCISION downto 1))+signed(MULTS_2_14(43)(PERCISION) & MULTS_2_14(43)(PERCISION downto 1));
			MULTS_3_7(44)<=signed(MULTS_2_13(44)(PERCISION) & MULTS_2_13(44)(PERCISION downto 1))+signed(MULTS_2_14(44)(PERCISION) & MULTS_2_14(44)(PERCISION downto 1));
			MULTS_3_7(45)<=signed(MULTS_2_13(45)(PERCISION) & MULTS_2_13(45)(PERCISION downto 1))+signed(MULTS_2_14(45)(PERCISION) & MULTS_2_14(45)(PERCISION downto 1));
			MULTS_3_7(46)<=signed(MULTS_2_13(46)(PERCISION) & MULTS_2_13(46)(PERCISION downto 1))+signed(MULTS_2_14(46)(PERCISION) & MULTS_2_14(46)(PERCISION downto 1));
			MULTS_3_7(47)<=signed(MULTS_2_13(47)(PERCISION) & MULTS_2_13(47)(PERCISION downto 1))+signed(MULTS_2_14(47)(PERCISION) & MULTS_2_14(47)(PERCISION downto 1));
			MULTS_3_7(48)<=signed(MULTS_2_13(48)(PERCISION) & MULTS_2_13(48)(PERCISION downto 1))+signed(MULTS_2_14(48)(PERCISION) & MULTS_2_14(48)(PERCISION downto 1));
			MULTS_3_7(49)<=signed(MULTS_2_13(49)(PERCISION) & MULTS_2_13(49)(PERCISION downto 1))+signed(MULTS_2_14(49)(PERCISION) & MULTS_2_14(49)(PERCISION downto 1));
			MULTS_3_7(50)<=signed(MULTS_2_13(50)(PERCISION) & MULTS_2_13(50)(PERCISION downto 1))+signed(MULTS_2_14(50)(PERCISION) & MULTS_2_14(50)(PERCISION downto 1));
			MULTS_3_7(51)<=signed(MULTS_2_13(51)(PERCISION) & MULTS_2_13(51)(PERCISION downto 1))+signed(MULTS_2_14(51)(PERCISION) & MULTS_2_14(51)(PERCISION downto 1));
			MULTS_3_7(52)<=signed(MULTS_2_13(52)(PERCISION) & MULTS_2_13(52)(PERCISION downto 1))+signed(MULTS_2_14(52)(PERCISION) & MULTS_2_14(52)(PERCISION downto 1));
			MULTS_3_7(53)<=signed(MULTS_2_13(53)(PERCISION) & MULTS_2_13(53)(PERCISION downto 1))+signed(MULTS_2_14(53)(PERCISION) & MULTS_2_14(53)(PERCISION downto 1));
			MULTS_3_7(54)<=signed(MULTS_2_13(54)(PERCISION) & MULTS_2_13(54)(PERCISION downto 1))+signed(MULTS_2_14(54)(PERCISION) & MULTS_2_14(54)(PERCISION downto 1));
			MULTS_3_7(55)<=signed(MULTS_2_13(55)(PERCISION) & MULTS_2_13(55)(PERCISION downto 1))+signed(MULTS_2_14(55)(PERCISION) & MULTS_2_14(55)(PERCISION downto 1));
			MULTS_3_7(56)<=signed(MULTS_2_13(56)(PERCISION) & MULTS_2_13(56)(PERCISION downto 1))+signed(MULTS_2_14(56)(PERCISION) & MULTS_2_14(56)(PERCISION downto 1));
			MULTS_3_7(57)<=signed(MULTS_2_13(57)(PERCISION) & MULTS_2_13(57)(PERCISION downto 1))+signed(MULTS_2_14(57)(PERCISION) & MULTS_2_14(57)(PERCISION downto 1));
			MULTS_3_7(58)<=signed(MULTS_2_13(58)(PERCISION) & MULTS_2_13(58)(PERCISION downto 1))+signed(MULTS_2_14(58)(PERCISION) & MULTS_2_14(58)(PERCISION downto 1));
			MULTS_3_7(59)<=signed(MULTS_2_13(59)(PERCISION) & MULTS_2_13(59)(PERCISION downto 1))+signed(MULTS_2_14(59)(PERCISION) & MULTS_2_14(59)(PERCISION downto 1));
			MULTS_3_7(60)<=signed(MULTS_2_13(60)(PERCISION) & MULTS_2_13(60)(PERCISION downto 1))+signed(MULTS_2_14(60)(PERCISION) & MULTS_2_14(60)(PERCISION downto 1));
			MULTS_3_7(61)<=signed(MULTS_2_13(61)(PERCISION) & MULTS_2_13(61)(PERCISION downto 1))+signed(MULTS_2_14(61)(PERCISION) & MULTS_2_14(61)(PERCISION downto 1));
			MULTS_3_7(62)<=signed(MULTS_2_13(62)(PERCISION) & MULTS_2_13(62)(PERCISION downto 1))+signed(MULTS_2_14(62)(PERCISION) & MULTS_2_14(62)(PERCISION downto 1));
			MULTS_3_7(63)<=signed(MULTS_2_13(63)(PERCISION) & MULTS_2_13(63)(PERCISION downto 1))+signed(MULTS_2_14(63)(PERCISION) & MULTS_2_14(63)(PERCISION downto 1));
			MULTS_3_7(64)<=signed(MULTS_2_13(64)(PERCISION) & MULTS_2_13(64)(PERCISION downto 1))+signed(MULTS_2_14(64)(PERCISION) & MULTS_2_14(64)(PERCISION downto 1));
			MULTS_3_7(65)<=signed(MULTS_2_13(65)(PERCISION) & MULTS_2_13(65)(PERCISION downto 1))+signed(MULTS_2_14(65)(PERCISION) & MULTS_2_14(65)(PERCISION downto 1));
			MULTS_3_7(66)<=signed(MULTS_2_13(66)(PERCISION) & MULTS_2_13(66)(PERCISION downto 1))+signed(MULTS_2_14(66)(PERCISION) & MULTS_2_14(66)(PERCISION downto 1));
			MULTS_3_7(67)<=signed(MULTS_2_13(67)(PERCISION) & MULTS_2_13(67)(PERCISION downto 1))+signed(MULTS_2_14(67)(PERCISION) & MULTS_2_14(67)(PERCISION downto 1));
			MULTS_3_7(68)<=signed(MULTS_2_13(68)(PERCISION) & MULTS_2_13(68)(PERCISION downto 1))+signed(MULTS_2_14(68)(PERCISION) & MULTS_2_14(68)(PERCISION downto 1));
			MULTS_3_7(69)<=signed(MULTS_2_13(69)(PERCISION) & MULTS_2_13(69)(PERCISION downto 1))+signed(MULTS_2_14(69)(PERCISION) & MULTS_2_14(69)(PERCISION downto 1));
			MULTS_3_7(70)<=signed(MULTS_2_13(70)(PERCISION) & MULTS_2_13(70)(PERCISION downto 1))+signed(MULTS_2_14(70)(PERCISION) & MULTS_2_14(70)(PERCISION downto 1));
			MULTS_3_7(71)<=signed(MULTS_2_13(71)(PERCISION) & MULTS_2_13(71)(PERCISION downto 1))+signed(MULTS_2_14(71)(PERCISION) & MULTS_2_14(71)(PERCISION downto 1));
			MULTS_3_7(72)<=signed(MULTS_2_13(72)(PERCISION) & MULTS_2_13(72)(PERCISION downto 1))+signed(MULTS_2_14(72)(PERCISION) & MULTS_2_14(72)(PERCISION downto 1));
			MULTS_3_7(73)<=signed(MULTS_2_13(73)(PERCISION) & MULTS_2_13(73)(PERCISION downto 1))+signed(MULTS_2_14(73)(PERCISION) & MULTS_2_14(73)(PERCISION downto 1));
			MULTS_3_7(74)<=signed(MULTS_2_13(74)(PERCISION) & MULTS_2_13(74)(PERCISION downto 1))+signed(MULTS_2_14(74)(PERCISION) & MULTS_2_14(74)(PERCISION downto 1));
			MULTS_3_7(75)<=signed(MULTS_2_13(75)(PERCISION) & MULTS_2_13(75)(PERCISION downto 1))+signed(MULTS_2_14(75)(PERCISION) & MULTS_2_14(75)(PERCISION downto 1));
			MULTS_3_7(76)<=signed(MULTS_2_13(76)(PERCISION) & MULTS_2_13(76)(PERCISION downto 1))+signed(MULTS_2_14(76)(PERCISION) & MULTS_2_14(76)(PERCISION downto 1));
			MULTS_3_7(77)<=signed(MULTS_2_13(77)(PERCISION) & MULTS_2_13(77)(PERCISION downto 1))+signed(MULTS_2_14(77)(PERCISION) & MULTS_2_14(77)(PERCISION downto 1));
			MULTS_3_7(78)<=signed(MULTS_2_13(78)(PERCISION) & MULTS_2_13(78)(PERCISION downto 1))+signed(MULTS_2_14(78)(PERCISION) & MULTS_2_14(78)(PERCISION downto 1));
			MULTS_3_7(79)<=signed(MULTS_2_13(79)(PERCISION) & MULTS_2_13(79)(PERCISION downto 1))+signed(MULTS_2_14(79)(PERCISION) & MULTS_2_14(79)(PERCISION downto 1));
			MULTS_3_7(80)<=signed(MULTS_2_13(80)(PERCISION) & MULTS_2_13(80)(PERCISION downto 1))+signed(MULTS_2_14(80)(PERCISION) & MULTS_2_14(80)(PERCISION downto 1));
			MULTS_3_7(81)<=signed(MULTS_2_13(81)(PERCISION) & MULTS_2_13(81)(PERCISION downto 1))+signed(MULTS_2_14(81)(PERCISION) & MULTS_2_14(81)(PERCISION downto 1));
			MULTS_3_7(82)<=signed(MULTS_2_13(82)(PERCISION) & MULTS_2_13(82)(PERCISION downto 1))+signed(MULTS_2_14(82)(PERCISION) & MULTS_2_14(82)(PERCISION downto 1));
			MULTS_3_7(83)<=signed(MULTS_2_13(83)(PERCISION) & MULTS_2_13(83)(PERCISION downto 1))+signed(MULTS_2_14(83)(PERCISION) & MULTS_2_14(83)(PERCISION downto 1));

			MULTS_3_8(0)<=signed(MULTS_2_15(0)(PERCISION) & MULTS_2_15(0)(PERCISION downto 1))+signed(MULTS_2_16(0)(PERCISION) & MULTS_2_16(0)(PERCISION downto 1));
			MULTS_3_8(1)<=signed(MULTS_2_15(1)(PERCISION) & MULTS_2_15(1)(PERCISION downto 1))+signed(MULTS_2_16(1)(PERCISION) & MULTS_2_16(1)(PERCISION downto 1));
			MULTS_3_8(2)<=signed(MULTS_2_15(2)(PERCISION) & MULTS_2_15(2)(PERCISION downto 1))+signed(MULTS_2_16(2)(PERCISION) & MULTS_2_16(2)(PERCISION downto 1));
			MULTS_3_8(3)<=signed(MULTS_2_15(3)(PERCISION) & MULTS_2_15(3)(PERCISION downto 1))+signed(MULTS_2_16(3)(PERCISION) & MULTS_2_16(3)(PERCISION downto 1));
			MULTS_3_8(4)<=signed(MULTS_2_15(4)(PERCISION) & MULTS_2_15(4)(PERCISION downto 1))+signed(MULTS_2_16(4)(PERCISION) & MULTS_2_16(4)(PERCISION downto 1));
			MULTS_3_8(5)<=signed(MULTS_2_15(5)(PERCISION) & MULTS_2_15(5)(PERCISION downto 1))+signed(MULTS_2_16(5)(PERCISION) & MULTS_2_16(5)(PERCISION downto 1));
			MULTS_3_8(6)<=signed(MULTS_2_15(6)(PERCISION) & MULTS_2_15(6)(PERCISION downto 1))+signed(MULTS_2_16(6)(PERCISION) & MULTS_2_16(6)(PERCISION downto 1));
			MULTS_3_8(7)<=signed(MULTS_2_15(7)(PERCISION) & MULTS_2_15(7)(PERCISION downto 1))+signed(MULTS_2_16(7)(PERCISION) & MULTS_2_16(7)(PERCISION downto 1));
			MULTS_3_8(8)<=signed(MULTS_2_15(8)(PERCISION) & MULTS_2_15(8)(PERCISION downto 1))+signed(MULTS_2_16(8)(PERCISION) & MULTS_2_16(8)(PERCISION downto 1));
			MULTS_3_8(9)<=signed(MULTS_2_15(9)(PERCISION) & MULTS_2_15(9)(PERCISION downto 1))+signed(MULTS_2_16(9)(PERCISION) & MULTS_2_16(9)(PERCISION downto 1));
			MULTS_3_8(10)<=signed(MULTS_2_15(10)(PERCISION) & MULTS_2_15(10)(PERCISION downto 1))+signed(MULTS_2_16(10)(PERCISION) & MULTS_2_16(10)(PERCISION downto 1));
			MULTS_3_8(11)<=signed(MULTS_2_15(11)(PERCISION) & MULTS_2_15(11)(PERCISION downto 1))+signed(MULTS_2_16(11)(PERCISION) & MULTS_2_16(11)(PERCISION downto 1));
			MULTS_3_8(12)<=signed(MULTS_2_15(12)(PERCISION) & MULTS_2_15(12)(PERCISION downto 1))+signed(MULTS_2_16(12)(PERCISION) & MULTS_2_16(12)(PERCISION downto 1));
			MULTS_3_8(13)<=signed(MULTS_2_15(13)(PERCISION) & MULTS_2_15(13)(PERCISION downto 1))+signed(MULTS_2_16(13)(PERCISION) & MULTS_2_16(13)(PERCISION downto 1));
			MULTS_3_8(14)<=signed(MULTS_2_15(14)(PERCISION) & MULTS_2_15(14)(PERCISION downto 1))+signed(MULTS_2_16(14)(PERCISION) & MULTS_2_16(14)(PERCISION downto 1));
			MULTS_3_8(15)<=signed(MULTS_2_15(15)(PERCISION) & MULTS_2_15(15)(PERCISION downto 1))+signed(MULTS_2_16(15)(PERCISION) & MULTS_2_16(15)(PERCISION downto 1));
			MULTS_3_8(16)<=signed(MULTS_2_15(16)(PERCISION) & MULTS_2_15(16)(PERCISION downto 1))+signed(MULTS_2_16(16)(PERCISION) & MULTS_2_16(16)(PERCISION downto 1));
			MULTS_3_8(17)<=signed(MULTS_2_15(17)(PERCISION) & MULTS_2_15(17)(PERCISION downto 1))+signed(MULTS_2_16(17)(PERCISION) & MULTS_2_16(17)(PERCISION downto 1));
			MULTS_3_8(18)<=signed(MULTS_2_15(18)(PERCISION) & MULTS_2_15(18)(PERCISION downto 1))+signed(MULTS_2_16(18)(PERCISION) & MULTS_2_16(18)(PERCISION downto 1));
			MULTS_3_8(19)<=signed(MULTS_2_15(19)(PERCISION) & MULTS_2_15(19)(PERCISION downto 1))+signed(MULTS_2_16(19)(PERCISION) & MULTS_2_16(19)(PERCISION downto 1));
			MULTS_3_8(20)<=signed(MULTS_2_15(20)(PERCISION) & MULTS_2_15(20)(PERCISION downto 1))+signed(MULTS_2_16(20)(PERCISION) & MULTS_2_16(20)(PERCISION downto 1));
			MULTS_3_8(21)<=signed(MULTS_2_15(21)(PERCISION) & MULTS_2_15(21)(PERCISION downto 1))+signed(MULTS_2_16(21)(PERCISION) & MULTS_2_16(21)(PERCISION downto 1));
			MULTS_3_8(22)<=signed(MULTS_2_15(22)(PERCISION) & MULTS_2_15(22)(PERCISION downto 1))+signed(MULTS_2_16(22)(PERCISION) & MULTS_2_16(22)(PERCISION downto 1));
			MULTS_3_8(23)<=signed(MULTS_2_15(23)(PERCISION) & MULTS_2_15(23)(PERCISION downto 1))+signed(MULTS_2_16(23)(PERCISION) & MULTS_2_16(23)(PERCISION downto 1));
			MULTS_3_8(24)<=signed(MULTS_2_15(24)(PERCISION) & MULTS_2_15(24)(PERCISION downto 1))+signed(MULTS_2_16(24)(PERCISION) & MULTS_2_16(24)(PERCISION downto 1));
			MULTS_3_8(25)<=signed(MULTS_2_15(25)(PERCISION) & MULTS_2_15(25)(PERCISION downto 1))+signed(MULTS_2_16(25)(PERCISION) & MULTS_2_16(25)(PERCISION downto 1));
			MULTS_3_8(26)<=signed(MULTS_2_15(26)(PERCISION) & MULTS_2_15(26)(PERCISION downto 1))+signed(MULTS_2_16(26)(PERCISION) & MULTS_2_16(26)(PERCISION downto 1));
			MULTS_3_8(27)<=signed(MULTS_2_15(27)(PERCISION) & MULTS_2_15(27)(PERCISION downto 1))+signed(MULTS_2_16(27)(PERCISION) & MULTS_2_16(27)(PERCISION downto 1));
			MULTS_3_8(28)<=signed(MULTS_2_15(28)(PERCISION) & MULTS_2_15(28)(PERCISION downto 1))+signed(MULTS_2_16(28)(PERCISION) & MULTS_2_16(28)(PERCISION downto 1));
			MULTS_3_8(29)<=signed(MULTS_2_15(29)(PERCISION) & MULTS_2_15(29)(PERCISION downto 1))+signed(MULTS_2_16(29)(PERCISION) & MULTS_2_16(29)(PERCISION downto 1));
			MULTS_3_8(30)<=signed(MULTS_2_15(30)(PERCISION) & MULTS_2_15(30)(PERCISION downto 1))+signed(MULTS_2_16(30)(PERCISION) & MULTS_2_16(30)(PERCISION downto 1));
			MULTS_3_8(31)<=signed(MULTS_2_15(31)(PERCISION) & MULTS_2_15(31)(PERCISION downto 1))+signed(MULTS_2_16(31)(PERCISION) & MULTS_2_16(31)(PERCISION downto 1));
			MULTS_3_8(32)<=signed(MULTS_2_15(32)(PERCISION) & MULTS_2_15(32)(PERCISION downto 1))+signed(MULTS_2_16(32)(PERCISION) & MULTS_2_16(32)(PERCISION downto 1));
			MULTS_3_8(33)<=signed(MULTS_2_15(33)(PERCISION) & MULTS_2_15(33)(PERCISION downto 1))+signed(MULTS_2_16(33)(PERCISION) & MULTS_2_16(33)(PERCISION downto 1));
			MULTS_3_8(34)<=signed(MULTS_2_15(34)(PERCISION) & MULTS_2_15(34)(PERCISION downto 1))+signed(MULTS_2_16(34)(PERCISION) & MULTS_2_16(34)(PERCISION downto 1));
			MULTS_3_8(35)<=signed(MULTS_2_15(35)(PERCISION) & MULTS_2_15(35)(PERCISION downto 1))+signed(MULTS_2_16(35)(PERCISION) & MULTS_2_16(35)(PERCISION downto 1));
			MULTS_3_8(36)<=signed(MULTS_2_15(36)(PERCISION) & MULTS_2_15(36)(PERCISION downto 1))+signed(MULTS_2_16(36)(PERCISION) & MULTS_2_16(36)(PERCISION downto 1));
			MULTS_3_8(37)<=signed(MULTS_2_15(37)(PERCISION) & MULTS_2_15(37)(PERCISION downto 1))+signed(MULTS_2_16(37)(PERCISION) & MULTS_2_16(37)(PERCISION downto 1));
			MULTS_3_8(38)<=signed(MULTS_2_15(38)(PERCISION) & MULTS_2_15(38)(PERCISION downto 1))+signed(MULTS_2_16(38)(PERCISION) & MULTS_2_16(38)(PERCISION downto 1));
			MULTS_3_8(39)<=signed(MULTS_2_15(39)(PERCISION) & MULTS_2_15(39)(PERCISION downto 1))+signed(MULTS_2_16(39)(PERCISION) & MULTS_2_16(39)(PERCISION downto 1));
			MULTS_3_8(40)<=signed(MULTS_2_15(40)(PERCISION) & MULTS_2_15(40)(PERCISION downto 1))+signed(MULTS_2_16(40)(PERCISION) & MULTS_2_16(40)(PERCISION downto 1));
			MULTS_3_8(41)<=signed(MULTS_2_15(41)(PERCISION) & MULTS_2_15(41)(PERCISION downto 1))+signed(MULTS_2_16(41)(PERCISION) & MULTS_2_16(41)(PERCISION downto 1));
			MULTS_3_8(42)<=signed(MULTS_2_15(42)(PERCISION) & MULTS_2_15(42)(PERCISION downto 1))+signed(MULTS_2_16(42)(PERCISION) & MULTS_2_16(42)(PERCISION downto 1));
			MULTS_3_8(43)<=signed(MULTS_2_15(43)(PERCISION) & MULTS_2_15(43)(PERCISION downto 1))+signed(MULTS_2_16(43)(PERCISION) & MULTS_2_16(43)(PERCISION downto 1));
			MULTS_3_8(44)<=signed(MULTS_2_15(44)(PERCISION) & MULTS_2_15(44)(PERCISION downto 1))+signed(MULTS_2_16(44)(PERCISION) & MULTS_2_16(44)(PERCISION downto 1));
			MULTS_3_8(45)<=signed(MULTS_2_15(45)(PERCISION) & MULTS_2_15(45)(PERCISION downto 1))+signed(MULTS_2_16(45)(PERCISION) & MULTS_2_16(45)(PERCISION downto 1));
			MULTS_3_8(46)<=signed(MULTS_2_15(46)(PERCISION) & MULTS_2_15(46)(PERCISION downto 1))+signed(MULTS_2_16(46)(PERCISION) & MULTS_2_16(46)(PERCISION downto 1));
			MULTS_3_8(47)<=signed(MULTS_2_15(47)(PERCISION) & MULTS_2_15(47)(PERCISION downto 1))+signed(MULTS_2_16(47)(PERCISION) & MULTS_2_16(47)(PERCISION downto 1));
			MULTS_3_8(48)<=signed(MULTS_2_15(48)(PERCISION) & MULTS_2_15(48)(PERCISION downto 1))+signed(MULTS_2_16(48)(PERCISION) & MULTS_2_16(48)(PERCISION downto 1));
			MULTS_3_8(49)<=signed(MULTS_2_15(49)(PERCISION) & MULTS_2_15(49)(PERCISION downto 1))+signed(MULTS_2_16(49)(PERCISION) & MULTS_2_16(49)(PERCISION downto 1));
			MULTS_3_8(50)<=signed(MULTS_2_15(50)(PERCISION) & MULTS_2_15(50)(PERCISION downto 1))+signed(MULTS_2_16(50)(PERCISION) & MULTS_2_16(50)(PERCISION downto 1));
			MULTS_3_8(51)<=signed(MULTS_2_15(51)(PERCISION) & MULTS_2_15(51)(PERCISION downto 1))+signed(MULTS_2_16(51)(PERCISION) & MULTS_2_16(51)(PERCISION downto 1));
			MULTS_3_8(52)<=signed(MULTS_2_15(52)(PERCISION) & MULTS_2_15(52)(PERCISION downto 1))+signed(MULTS_2_16(52)(PERCISION) & MULTS_2_16(52)(PERCISION downto 1));
			MULTS_3_8(53)<=signed(MULTS_2_15(53)(PERCISION) & MULTS_2_15(53)(PERCISION downto 1))+signed(MULTS_2_16(53)(PERCISION) & MULTS_2_16(53)(PERCISION downto 1));
			MULTS_3_8(54)<=signed(MULTS_2_15(54)(PERCISION) & MULTS_2_15(54)(PERCISION downto 1))+signed(MULTS_2_16(54)(PERCISION) & MULTS_2_16(54)(PERCISION downto 1));
			MULTS_3_8(55)<=signed(MULTS_2_15(55)(PERCISION) & MULTS_2_15(55)(PERCISION downto 1))+signed(MULTS_2_16(55)(PERCISION) & MULTS_2_16(55)(PERCISION downto 1));
			MULTS_3_8(56)<=signed(MULTS_2_15(56)(PERCISION) & MULTS_2_15(56)(PERCISION downto 1))+signed(MULTS_2_16(56)(PERCISION) & MULTS_2_16(56)(PERCISION downto 1));
			MULTS_3_8(57)<=signed(MULTS_2_15(57)(PERCISION) & MULTS_2_15(57)(PERCISION downto 1))+signed(MULTS_2_16(57)(PERCISION) & MULTS_2_16(57)(PERCISION downto 1));
			MULTS_3_8(58)<=signed(MULTS_2_15(58)(PERCISION) & MULTS_2_15(58)(PERCISION downto 1))+signed(MULTS_2_16(58)(PERCISION) & MULTS_2_16(58)(PERCISION downto 1));
			MULTS_3_8(59)<=signed(MULTS_2_15(59)(PERCISION) & MULTS_2_15(59)(PERCISION downto 1))+signed(MULTS_2_16(59)(PERCISION) & MULTS_2_16(59)(PERCISION downto 1));
			MULTS_3_8(60)<=signed(MULTS_2_15(60)(PERCISION) & MULTS_2_15(60)(PERCISION downto 1))+signed(MULTS_2_16(60)(PERCISION) & MULTS_2_16(60)(PERCISION downto 1));
			MULTS_3_8(61)<=signed(MULTS_2_15(61)(PERCISION) & MULTS_2_15(61)(PERCISION downto 1))+signed(MULTS_2_16(61)(PERCISION) & MULTS_2_16(61)(PERCISION downto 1));
			MULTS_3_8(62)<=signed(MULTS_2_15(62)(PERCISION) & MULTS_2_15(62)(PERCISION downto 1))+signed(MULTS_2_16(62)(PERCISION) & MULTS_2_16(62)(PERCISION downto 1));
			MULTS_3_8(63)<=signed(MULTS_2_15(63)(PERCISION) & MULTS_2_15(63)(PERCISION downto 1))+signed(MULTS_2_16(63)(PERCISION) & MULTS_2_16(63)(PERCISION downto 1));
			MULTS_3_8(64)<=signed(MULTS_2_15(64)(PERCISION) & MULTS_2_15(64)(PERCISION downto 1))+signed(MULTS_2_16(64)(PERCISION) & MULTS_2_16(64)(PERCISION downto 1));
			MULTS_3_8(65)<=signed(MULTS_2_15(65)(PERCISION) & MULTS_2_15(65)(PERCISION downto 1))+signed(MULTS_2_16(65)(PERCISION) & MULTS_2_16(65)(PERCISION downto 1));
			MULTS_3_8(66)<=signed(MULTS_2_15(66)(PERCISION) & MULTS_2_15(66)(PERCISION downto 1))+signed(MULTS_2_16(66)(PERCISION) & MULTS_2_16(66)(PERCISION downto 1));
			MULTS_3_8(67)<=signed(MULTS_2_15(67)(PERCISION) & MULTS_2_15(67)(PERCISION downto 1))+signed(MULTS_2_16(67)(PERCISION) & MULTS_2_16(67)(PERCISION downto 1));
			MULTS_3_8(68)<=signed(MULTS_2_15(68)(PERCISION) & MULTS_2_15(68)(PERCISION downto 1))+signed(MULTS_2_16(68)(PERCISION) & MULTS_2_16(68)(PERCISION downto 1));
			MULTS_3_8(69)<=signed(MULTS_2_15(69)(PERCISION) & MULTS_2_15(69)(PERCISION downto 1))+signed(MULTS_2_16(69)(PERCISION) & MULTS_2_16(69)(PERCISION downto 1));
			MULTS_3_8(70)<=signed(MULTS_2_15(70)(PERCISION) & MULTS_2_15(70)(PERCISION downto 1))+signed(MULTS_2_16(70)(PERCISION) & MULTS_2_16(70)(PERCISION downto 1));
			MULTS_3_8(71)<=signed(MULTS_2_15(71)(PERCISION) & MULTS_2_15(71)(PERCISION downto 1))+signed(MULTS_2_16(71)(PERCISION) & MULTS_2_16(71)(PERCISION downto 1));
			MULTS_3_8(72)<=signed(MULTS_2_15(72)(PERCISION) & MULTS_2_15(72)(PERCISION downto 1))+signed(MULTS_2_16(72)(PERCISION) & MULTS_2_16(72)(PERCISION downto 1));
			MULTS_3_8(73)<=signed(MULTS_2_15(73)(PERCISION) & MULTS_2_15(73)(PERCISION downto 1))+signed(MULTS_2_16(73)(PERCISION) & MULTS_2_16(73)(PERCISION downto 1));
			MULTS_3_8(74)<=signed(MULTS_2_15(74)(PERCISION) & MULTS_2_15(74)(PERCISION downto 1))+signed(MULTS_2_16(74)(PERCISION) & MULTS_2_16(74)(PERCISION downto 1));
			MULTS_3_8(75)<=signed(MULTS_2_15(75)(PERCISION) & MULTS_2_15(75)(PERCISION downto 1))+signed(MULTS_2_16(75)(PERCISION) & MULTS_2_16(75)(PERCISION downto 1));
			MULTS_3_8(76)<=signed(MULTS_2_15(76)(PERCISION) & MULTS_2_15(76)(PERCISION downto 1))+signed(MULTS_2_16(76)(PERCISION) & MULTS_2_16(76)(PERCISION downto 1));
			MULTS_3_8(77)<=signed(MULTS_2_15(77)(PERCISION) & MULTS_2_15(77)(PERCISION downto 1))+signed(MULTS_2_16(77)(PERCISION) & MULTS_2_16(77)(PERCISION downto 1));
			MULTS_3_8(78)<=signed(MULTS_2_15(78)(PERCISION) & MULTS_2_15(78)(PERCISION downto 1))+signed(MULTS_2_16(78)(PERCISION) & MULTS_2_16(78)(PERCISION downto 1));
			MULTS_3_8(79)<=signed(MULTS_2_15(79)(PERCISION) & MULTS_2_15(79)(PERCISION downto 1))+signed(MULTS_2_16(79)(PERCISION) & MULTS_2_16(79)(PERCISION downto 1));
			MULTS_3_8(80)<=signed(MULTS_2_15(80)(PERCISION) & MULTS_2_15(80)(PERCISION downto 1))+signed(MULTS_2_16(80)(PERCISION) & MULTS_2_16(80)(PERCISION downto 1));
			MULTS_3_8(81)<=signed(MULTS_2_15(81)(PERCISION) & MULTS_2_15(81)(PERCISION downto 1))+signed(MULTS_2_16(81)(PERCISION) & MULTS_2_16(81)(PERCISION downto 1));
			MULTS_3_8(82)<=signed(MULTS_2_15(82)(PERCISION) & MULTS_2_15(82)(PERCISION downto 1))+signed(MULTS_2_16(82)(PERCISION) & MULTS_2_16(82)(PERCISION downto 1));
			MULTS_3_8(83)<=signed(MULTS_2_15(83)(PERCISION) & MULTS_2_15(83)(PERCISION downto 1))+signed(MULTS_2_16(83)(PERCISION) & MULTS_2_16(83)(PERCISION downto 1));



                         EN_SUM_MULT_4<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_4 = '1' then
			------------------------------------STAGE-4--------------------------------------
			MULTS_4_1(0)<=signed(MULTS_3_1(0));
			MULTS_4_1(1)<=signed(MULTS_3_1(1));
			MULTS_4_1(2)<=signed(MULTS_3_1(2));
			MULTS_4_1(3)<=signed(MULTS_3_1(3));
			MULTS_4_1(4)<=signed(MULTS_3_1(4));
			MULTS_4_1(5)<=signed(MULTS_3_1(5));
			MULTS_4_1(6)<=signed(MULTS_3_1(6));
			MULTS_4_1(7)<=signed(MULTS_3_1(7));
			MULTS_4_1(8)<=signed(MULTS_3_1(8));
			MULTS_4_1(9)<=signed(MULTS_3_1(9));
			MULTS_4_1(10)<=signed(MULTS_3_1(10));
			MULTS_4_1(11)<=signed(MULTS_3_1(11));
			MULTS_4_1(12)<=signed(MULTS_3_1(12));
			MULTS_4_1(13)<=signed(MULTS_3_1(13));
			MULTS_4_1(14)<=signed(MULTS_3_1(14));
			MULTS_4_1(15)<=signed(MULTS_3_1(15));
			MULTS_4_1(16)<=signed(MULTS_3_1(16));
			MULTS_4_1(17)<=signed(MULTS_3_1(17));
			MULTS_4_1(18)<=signed(MULTS_3_1(18));
			MULTS_4_1(19)<=signed(MULTS_3_1(19));
			MULTS_4_1(20)<=signed(MULTS_3_1(20));
			MULTS_4_1(21)<=signed(MULTS_3_1(21));
			MULTS_4_1(22)<=signed(MULTS_3_1(22));
			MULTS_4_1(23)<=signed(MULTS_3_1(23));
			MULTS_4_1(24)<=signed(MULTS_3_1(24));
			MULTS_4_1(25)<=signed(MULTS_3_1(25));
			MULTS_4_1(26)<=signed(MULTS_3_1(26));
			MULTS_4_1(27)<=signed(MULTS_3_1(27));
			MULTS_4_1(28)<=signed(MULTS_3_1(28));
			MULTS_4_1(29)<=signed(MULTS_3_1(29));
			MULTS_4_1(30)<=signed(MULTS_3_1(30));
			MULTS_4_1(31)<=signed(MULTS_3_1(31));
			MULTS_4_1(32)<=signed(MULTS_3_1(32));
			MULTS_4_1(33)<=signed(MULTS_3_1(33));
			MULTS_4_1(34)<=signed(MULTS_3_1(34));
			MULTS_4_1(35)<=signed(MULTS_3_1(35));
			MULTS_4_1(36)<=signed(MULTS_3_1(36));
			MULTS_4_1(37)<=signed(MULTS_3_1(37));
			MULTS_4_1(38)<=signed(MULTS_3_1(38));
			MULTS_4_1(39)<=signed(MULTS_3_1(39));
			MULTS_4_1(40)<=signed(MULTS_3_1(40));
			MULTS_4_1(41)<=signed(MULTS_3_1(41));
			MULTS_4_1(42)<=signed(MULTS_3_1(42));
			MULTS_4_1(43)<=signed(MULTS_3_1(43));
			MULTS_4_1(44)<=signed(MULTS_3_1(44));
			MULTS_4_1(45)<=signed(MULTS_3_1(45));
			MULTS_4_1(46)<=signed(MULTS_3_1(46));
			MULTS_4_1(47)<=signed(MULTS_3_1(47));
			MULTS_4_1(48)<=signed(MULTS_3_1(48));
			MULTS_4_1(49)<=signed(MULTS_3_1(49));
			MULTS_4_1(50)<=signed(MULTS_3_1(50));
			MULTS_4_1(51)<=signed(MULTS_3_1(51));
			MULTS_4_1(52)<=signed(MULTS_3_1(52));
			MULTS_4_1(53)<=signed(MULTS_3_1(53));
			MULTS_4_1(54)<=signed(MULTS_3_1(54));
			MULTS_4_1(55)<=signed(MULTS_3_1(55));
			MULTS_4_1(56)<=signed(MULTS_3_1(56));
			MULTS_4_1(57)<=signed(MULTS_3_1(57));
			MULTS_4_1(58)<=signed(MULTS_3_1(58));
			MULTS_4_1(59)<=signed(MULTS_3_1(59));
			MULTS_4_1(60)<=signed(MULTS_3_1(60));
			MULTS_4_1(61)<=signed(MULTS_3_1(61));
			MULTS_4_1(62)<=signed(MULTS_3_1(62));
			MULTS_4_1(63)<=signed(MULTS_3_1(63));
			MULTS_4_1(64)<=signed(MULTS_3_1(64));
			MULTS_4_1(65)<=signed(MULTS_3_1(65));
			MULTS_4_1(66)<=signed(MULTS_3_1(66));
			MULTS_4_1(67)<=signed(MULTS_3_1(67));
			MULTS_4_1(68)<=signed(MULTS_3_1(68));
			MULTS_4_1(69)<=signed(MULTS_3_1(69));
			MULTS_4_1(70)<=signed(MULTS_3_1(70));
			MULTS_4_1(71)<=signed(MULTS_3_1(71));
			MULTS_4_1(72)<=signed(MULTS_3_1(72));
			MULTS_4_1(73)<=signed(MULTS_3_1(73));
			MULTS_4_1(74)<=signed(MULTS_3_1(74));
			MULTS_4_1(75)<=signed(MULTS_3_1(75));
			MULTS_4_1(76)<=signed(MULTS_3_1(76));
			MULTS_4_1(77)<=signed(MULTS_3_1(77));
			MULTS_4_1(78)<=signed(MULTS_3_1(78));
			MULTS_4_1(79)<=signed(MULTS_3_1(79));
			MULTS_4_1(80)<=signed(MULTS_3_1(80));
			MULTS_4_1(81)<=signed(MULTS_3_1(81));
			MULTS_4_1(82)<=signed(MULTS_3_1(82));
			MULTS_4_1(83)<=signed(MULTS_3_1(83));

			MULTS_4_2(0)<=signed(MULTS_3_2(0)(PERCISION) & MULTS_3_2(0)(PERCISION downto 1))+signed(MULTS_3_3(0)(PERCISION) & MULTS_3_3(0)(PERCISION downto 1));
			MULTS_4_2(1)<=signed(MULTS_3_2(1)(PERCISION) & MULTS_3_2(1)(PERCISION downto 1))+signed(MULTS_3_3(1)(PERCISION) & MULTS_3_3(1)(PERCISION downto 1));
			MULTS_4_2(2)<=signed(MULTS_3_2(2)(PERCISION) & MULTS_3_2(2)(PERCISION downto 1))+signed(MULTS_3_3(2)(PERCISION) & MULTS_3_3(2)(PERCISION downto 1));
			MULTS_4_2(3)<=signed(MULTS_3_2(3)(PERCISION) & MULTS_3_2(3)(PERCISION downto 1))+signed(MULTS_3_3(3)(PERCISION) & MULTS_3_3(3)(PERCISION downto 1));
			MULTS_4_2(4)<=signed(MULTS_3_2(4)(PERCISION) & MULTS_3_2(4)(PERCISION downto 1))+signed(MULTS_3_3(4)(PERCISION) & MULTS_3_3(4)(PERCISION downto 1));
			MULTS_4_2(5)<=signed(MULTS_3_2(5)(PERCISION) & MULTS_3_2(5)(PERCISION downto 1))+signed(MULTS_3_3(5)(PERCISION) & MULTS_3_3(5)(PERCISION downto 1));
			MULTS_4_2(6)<=signed(MULTS_3_2(6)(PERCISION) & MULTS_3_2(6)(PERCISION downto 1))+signed(MULTS_3_3(6)(PERCISION) & MULTS_3_3(6)(PERCISION downto 1));
			MULTS_4_2(7)<=signed(MULTS_3_2(7)(PERCISION) & MULTS_3_2(7)(PERCISION downto 1))+signed(MULTS_3_3(7)(PERCISION) & MULTS_3_3(7)(PERCISION downto 1));
			MULTS_4_2(8)<=signed(MULTS_3_2(8)(PERCISION) & MULTS_3_2(8)(PERCISION downto 1))+signed(MULTS_3_3(8)(PERCISION) & MULTS_3_3(8)(PERCISION downto 1));
			MULTS_4_2(9)<=signed(MULTS_3_2(9)(PERCISION) & MULTS_3_2(9)(PERCISION downto 1))+signed(MULTS_3_3(9)(PERCISION) & MULTS_3_3(9)(PERCISION downto 1));
			MULTS_4_2(10)<=signed(MULTS_3_2(10)(PERCISION) & MULTS_3_2(10)(PERCISION downto 1))+signed(MULTS_3_3(10)(PERCISION) & MULTS_3_3(10)(PERCISION downto 1));
			MULTS_4_2(11)<=signed(MULTS_3_2(11)(PERCISION) & MULTS_3_2(11)(PERCISION downto 1))+signed(MULTS_3_3(11)(PERCISION) & MULTS_3_3(11)(PERCISION downto 1));
			MULTS_4_2(12)<=signed(MULTS_3_2(12)(PERCISION) & MULTS_3_2(12)(PERCISION downto 1))+signed(MULTS_3_3(12)(PERCISION) & MULTS_3_3(12)(PERCISION downto 1));
			MULTS_4_2(13)<=signed(MULTS_3_2(13)(PERCISION) & MULTS_3_2(13)(PERCISION downto 1))+signed(MULTS_3_3(13)(PERCISION) & MULTS_3_3(13)(PERCISION downto 1));
			MULTS_4_2(14)<=signed(MULTS_3_2(14)(PERCISION) & MULTS_3_2(14)(PERCISION downto 1))+signed(MULTS_3_3(14)(PERCISION) & MULTS_3_3(14)(PERCISION downto 1));
			MULTS_4_2(15)<=signed(MULTS_3_2(15)(PERCISION) & MULTS_3_2(15)(PERCISION downto 1))+signed(MULTS_3_3(15)(PERCISION) & MULTS_3_3(15)(PERCISION downto 1));
			MULTS_4_2(16)<=signed(MULTS_3_2(16)(PERCISION) & MULTS_3_2(16)(PERCISION downto 1))+signed(MULTS_3_3(16)(PERCISION) & MULTS_3_3(16)(PERCISION downto 1));
			MULTS_4_2(17)<=signed(MULTS_3_2(17)(PERCISION) & MULTS_3_2(17)(PERCISION downto 1))+signed(MULTS_3_3(17)(PERCISION) & MULTS_3_3(17)(PERCISION downto 1));
			MULTS_4_2(18)<=signed(MULTS_3_2(18)(PERCISION) & MULTS_3_2(18)(PERCISION downto 1))+signed(MULTS_3_3(18)(PERCISION) & MULTS_3_3(18)(PERCISION downto 1));
			MULTS_4_2(19)<=signed(MULTS_3_2(19)(PERCISION) & MULTS_3_2(19)(PERCISION downto 1))+signed(MULTS_3_3(19)(PERCISION) & MULTS_3_3(19)(PERCISION downto 1));
			MULTS_4_2(20)<=signed(MULTS_3_2(20)(PERCISION) & MULTS_3_2(20)(PERCISION downto 1))+signed(MULTS_3_3(20)(PERCISION) & MULTS_3_3(20)(PERCISION downto 1));
			MULTS_4_2(21)<=signed(MULTS_3_2(21)(PERCISION) & MULTS_3_2(21)(PERCISION downto 1))+signed(MULTS_3_3(21)(PERCISION) & MULTS_3_3(21)(PERCISION downto 1));
			MULTS_4_2(22)<=signed(MULTS_3_2(22)(PERCISION) & MULTS_3_2(22)(PERCISION downto 1))+signed(MULTS_3_3(22)(PERCISION) & MULTS_3_3(22)(PERCISION downto 1));
			MULTS_4_2(23)<=signed(MULTS_3_2(23)(PERCISION) & MULTS_3_2(23)(PERCISION downto 1))+signed(MULTS_3_3(23)(PERCISION) & MULTS_3_3(23)(PERCISION downto 1));
			MULTS_4_2(24)<=signed(MULTS_3_2(24)(PERCISION) & MULTS_3_2(24)(PERCISION downto 1))+signed(MULTS_3_3(24)(PERCISION) & MULTS_3_3(24)(PERCISION downto 1));
			MULTS_4_2(25)<=signed(MULTS_3_2(25)(PERCISION) & MULTS_3_2(25)(PERCISION downto 1))+signed(MULTS_3_3(25)(PERCISION) & MULTS_3_3(25)(PERCISION downto 1));
			MULTS_4_2(26)<=signed(MULTS_3_2(26)(PERCISION) & MULTS_3_2(26)(PERCISION downto 1))+signed(MULTS_3_3(26)(PERCISION) & MULTS_3_3(26)(PERCISION downto 1));
			MULTS_4_2(27)<=signed(MULTS_3_2(27)(PERCISION) & MULTS_3_2(27)(PERCISION downto 1))+signed(MULTS_3_3(27)(PERCISION) & MULTS_3_3(27)(PERCISION downto 1));
			MULTS_4_2(28)<=signed(MULTS_3_2(28)(PERCISION) & MULTS_3_2(28)(PERCISION downto 1))+signed(MULTS_3_3(28)(PERCISION) & MULTS_3_3(28)(PERCISION downto 1));
			MULTS_4_2(29)<=signed(MULTS_3_2(29)(PERCISION) & MULTS_3_2(29)(PERCISION downto 1))+signed(MULTS_3_3(29)(PERCISION) & MULTS_3_3(29)(PERCISION downto 1));
			MULTS_4_2(30)<=signed(MULTS_3_2(30)(PERCISION) & MULTS_3_2(30)(PERCISION downto 1))+signed(MULTS_3_3(30)(PERCISION) & MULTS_3_3(30)(PERCISION downto 1));
			MULTS_4_2(31)<=signed(MULTS_3_2(31)(PERCISION) & MULTS_3_2(31)(PERCISION downto 1))+signed(MULTS_3_3(31)(PERCISION) & MULTS_3_3(31)(PERCISION downto 1));
			MULTS_4_2(32)<=signed(MULTS_3_2(32)(PERCISION) & MULTS_3_2(32)(PERCISION downto 1))+signed(MULTS_3_3(32)(PERCISION) & MULTS_3_3(32)(PERCISION downto 1));
			MULTS_4_2(33)<=signed(MULTS_3_2(33)(PERCISION) & MULTS_3_2(33)(PERCISION downto 1))+signed(MULTS_3_3(33)(PERCISION) & MULTS_3_3(33)(PERCISION downto 1));
			MULTS_4_2(34)<=signed(MULTS_3_2(34)(PERCISION) & MULTS_3_2(34)(PERCISION downto 1))+signed(MULTS_3_3(34)(PERCISION) & MULTS_3_3(34)(PERCISION downto 1));
			MULTS_4_2(35)<=signed(MULTS_3_2(35)(PERCISION) & MULTS_3_2(35)(PERCISION downto 1))+signed(MULTS_3_3(35)(PERCISION) & MULTS_3_3(35)(PERCISION downto 1));
			MULTS_4_2(36)<=signed(MULTS_3_2(36)(PERCISION) & MULTS_3_2(36)(PERCISION downto 1))+signed(MULTS_3_3(36)(PERCISION) & MULTS_3_3(36)(PERCISION downto 1));
			MULTS_4_2(37)<=signed(MULTS_3_2(37)(PERCISION) & MULTS_3_2(37)(PERCISION downto 1))+signed(MULTS_3_3(37)(PERCISION) & MULTS_3_3(37)(PERCISION downto 1));
			MULTS_4_2(38)<=signed(MULTS_3_2(38)(PERCISION) & MULTS_3_2(38)(PERCISION downto 1))+signed(MULTS_3_3(38)(PERCISION) & MULTS_3_3(38)(PERCISION downto 1));
			MULTS_4_2(39)<=signed(MULTS_3_2(39)(PERCISION) & MULTS_3_2(39)(PERCISION downto 1))+signed(MULTS_3_3(39)(PERCISION) & MULTS_3_3(39)(PERCISION downto 1));
			MULTS_4_2(40)<=signed(MULTS_3_2(40)(PERCISION) & MULTS_3_2(40)(PERCISION downto 1))+signed(MULTS_3_3(40)(PERCISION) & MULTS_3_3(40)(PERCISION downto 1));
			MULTS_4_2(41)<=signed(MULTS_3_2(41)(PERCISION) & MULTS_3_2(41)(PERCISION downto 1))+signed(MULTS_3_3(41)(PERCISION) & MULTS_3_3(41)(PERCISION downto 1));
			MULTS_4_2(42)<=signed(MULTS_3_2(42)(PERCISION) & MULTS_3_2(42)(PERCISION downto 1))+signed(MULTS_3_3(42)(PERCISION) & MULTS_3_3(42)(PERCISION downto 1));
			MULTS_4_2(43)<=signed(MULTS_3_2(43)(PERCISION) & MULTS_3_2(43)(PERCISION downto 1))+signed(MULTS_3_3(43)(PERCISION) & MULTS_3_3(43)(PERCISION downto 1));
			MULTS_4_2(44)<=signed(MULTS_3_2(44)(PERCISION) & MULTS_3_2(44)(PERCISION downto 1))+signed(MULTS_3_3(44)(PERCISION) & MULTS_3_3(44)(PERCISION downto 1));
			MULTS_4_2(45)<=signed(MULTS_3_2(45)(PERCISION) & MULTS_3_2(45)(PERCISION downto 1))+signed(MULTS_3_3(45)(PERCISION) & MULTS_3_3(45)(PERCISION downto 1));
			MULTS_4_2(46)<=signed(MULTS_3_2(46)(PERCISION) & MULTS_3_2(46)(PERCISION downto 1))+signed(MULTS_3_3(46)(PERCISION) & MULTS_3_3(46)(PERCISION downto 1));
			MULTS_4_2(47)<=signed(MULTS_3_2(47)(PERCISION) & MULTS_3_2(47)(PERCISION downto 1))+signed(MULTS_3_3(47)(PERCISION) & MULTS_3_3(47)(PERCISION downto 1));
			MULTS_4_2(48)<=signed(MULTS_3_2(48)(PERCISION) & MULTS_3_2(48)(PERCISION downto 1))+signed(MULTS_3_3(48)(PERCISION) & MULTS_3_3(48)(PERCISION downto 1));
			MULTS_4_2(49)<=signed(MULTS_3_2(49)(PERCISION) & MULTS_3_2(49)(PERCISION downto 1))+signed(MULTS_3_3(49)(PERCISION) & MULTS_3_3(49)(PERCISION downto 1));
			MULTS_4_2(50)<=signed(MULTS_3_2(50)(PERCISION) & MULTS_3_2(50)(PERCISION downto 1))+signed(MULTS_3_3(50)(PERCISION) & MULTS_3_3(50)(PERCISION downto 1));
			MULTS_4_2(51)<=signed(MULTS_3_2(51)(PERCISION) & MULTS_3_2(51)(PERCISION downto 1))+signed(MULTS_3_3(51)(PERCISION) & MULTS_3_3(51)(PERCISION downto 1));
			MULTS_4_2(52)<=signed(MULTS_3_2(52)(PERCISION) & MULTS_3_2(52)(PERCISION downto 1))+signed(MULTS_3_3(52)(PERCISION) & MULTS_3_3(52)(PERCISION downto 1));
			MULTS_4_2(53)<=signed(MULTS_3_2(53)(PERCISION) & MULTS_3_2(53)(PERCISION downto 1))+signed(MULTS_3_3(53)(PERCISION) & MULTS_3_3(53)(PERCISION downto 1));
			MULTS_4_2(54)<=signed(MULTS_3_2(54)(PERCISION) & MULTS_3_2(54)(PERCISION downto 1))+signed(MULTS_3_3(54)(PERCISION) & MULTS_3_3(54)(PERCISION downto 1));
			MULTS_4_2(55)<=signed(MULTS_3_2(55)(PERCISION) & MULTS_3_2(55)(PERCISION downto 1))+signed(MULTS_3_3(55)(PERCISION) & MULTS_3_3(55)(PERCISION downto 1));
			MULTS_4_2(56)<=signed(MULTS_3_2(56)(PERCISION) & MULTS_3_2(56)(PERCISION downto 1))+signed(MULTS_3_3(56)(PERCISION) & MULTS_3_3(56)(PERCISION downto 1));
			MULTS_4_2(57)<=signed(MULTS_3_2(57)(PERCISION) & MULTS_3_2(57)(PERCISION downto 1))+signed(MULTS_3_3(57)(PERCISION) & MULTS_3_3(57)(PERCISION downto 1));
			MULTS_4_2(58)<=signed(MULTS_3_2(58)(PERCISION) & MULTS_3_2(58)(PERCISION downto 1))+signed(MULTS_3_3(58)(PERCISION) & MULTS_3_3(58)(PERCISION downto 1));
			MULTS_4_2(59)<=signed(MULTS_3_2(59)(PERCISION) & MULTS_3_2(59)(PERCISION downto 1))+signed(MULTS_3_3(59)(PERCISION) & MULTS_3_3(59)(PERCISION downto 1));
			MULTS_4_2(60)<=signed(MULTS_3_2(60)(PERCISION) & MULTS_3_2(60)(PERCISION downto 1))+signed(MULTS_3_3(60)(PERCISION) & MULTS_3_3(60)(PERCISION downto 1));
			MULTS_4_2(61)<=signed(MULTS_3_2(61)(PERCISION) & MULTS_3_2(61)(PERCISION downto 1))+signed(MULTS_3_3(61)(PERCISION) & MULTS_3_3(61)(PERCISION downto 1));
			MULTS_4_2(62)<=signed(MULTS_3_2(62)(PERCISION) & MULTS_3_2(62)(PERCISION downto 1))+signed(MULTS_3_3(62)(PERCISION) & MULTS_3_3(62)(PERCISION downto 1));
			MULTS_4_2(63)<=signed(MULTS_3_2(63)(PERCISION) & MULTS_3_2(63)(PERCISION downto 1))+signed(MULTS_3_3(63)(PERCISION) & MULTS_3_3(63)(PERCISION downto 1));
			MULTS_4_2(64)<=signed(MULTS_3_2(64)(PERCISION) & MULTS_3_2(64)(PERCISION downto 1))+signed(MULTS_3_3(64)(PERCISION) & MULTS_3_3(64)(PERCISION downto 1));
			MULTS_4_2(65)<=signed(MULTS_3_2(65)(PERCISION) & MULTS_3_2(65)(PERCISION downto 1))+signed(MULTS_3_3(65)(PERCISION) & MULTS_3_3(65)(PERCISION downto 1));
			MULTS_4_2(66)<=signed(MULTS_3_2(66)(PERCISION) & MULTS_3_2(66)(PERCISION downto 1))+signed(MULTS_3_3(66)(PERCISION) & MULTS_3_3(66)(PERCISION downto 1));
			MULTS_4_2(67)<=signed(MULTS_3_2(67)(PERCISION) & MULTS_3_2(67)(PERCISION downto 1))+signed(MULTS_3_3(67)(PERCISION) & MULTS_3_3(67)(PERCISION downto 1));
			MULTS_4_2(68)<=signed(MULTS_3_2(68)(PERCISION) & MULTS_3_2(68)(PERCISION downto 1))+signed(MULTS_3_3(68)(PERCISION) & MULTS_3_3(68)(PERCISION downto 1));
			MULTS_4_2(69)<=signed(MULTS_3_2(69)(PERCISION) & MULTS_3_2(69)(PERCISION downto 1))+signed(MULTS_3_3(69)(PERCISION) & MULTS_3_3(69)(PERCISION downto 1));
			MULTS_4_2(70)<=signed(MULTS_3_2(70)(PERCISION) & MULTS_3_2(70)(PERCISION downto 1))+signed(MULTS_3_3(70)(PERCISION) & MULTS_3_3(70)(PERCISION downto 1));
			MULTS_4_2(71)<=signed(MULTS_3_2(71)(PERCISION) & MULTS_3_2(71)(PERCISION downto 1))+signed(MULTS_3_3(71)(PERCISION) & MULTS_3_3(71)(PERCISION downto 1));
			MULTS_4_2(72)<=signed(MULTS_3_2(72)(PERCISION) & MULTS_3_2(72)(PERCISION downto 1))+signed(MULTS_3_3(72)(PERCISION) & MULTS_3_3(72)(PERCISION downto 1));
			MULTS_4_2(73)<=signed(MULTS_3_2(73)(PERCISION) & MULTS_3_2(73)(PERCISION downto 1))+signed(MULTS_3_3(73)(PERCISION) & MULTS_3_3(73)(PERCISION downto 1));
			MULTS_4_2(74)<=signed(MULTS_3_2(74)(PERCISION) & MULTS_3_2(74)(PERCISION downto 1))+signed(MULTS_3_3(74)(PERCISION) & MULTS_3_3(74)(PERCISION downto 1));
			MULTS_4_2(75)<=signed(MULTS_3_2(75)(PERCISION) & MULTS_3_2(75)(PERCISION downto 1))+signed(MULTS_3_3(75)(PERCISION) & MULTS_3_3(75)(PERCISION downto 1));
			MULTS_4_2(76)<=signed(MULTS_3_2(76)(PERCISION) & MULTS_3_2(76)(PERCISION downto 1))+signed(MULTS_3_3(76)(PERCISION) & MULTS_3_3(76)(PERCISION downto 1));
			MULTS_4_2(77)<=signed(MULTS_3_2(77)(PERCISION) & MULTS_3_2(77)(PERCISION downto 1))+signed(MULTS_3_3(77)(PERCISION) & MULTS_3_3(77)(PERCISION downto 1));
			MULTS_4_2(78)<=signed(MULTS_3_2(78)(PERCISION) & MULTS_3_2(78)(PERCISION downto 1))+signed(MULTS_3_3(78)(PERCISION) & MULTS_3_3(78)(PERCISION downto 1));
			MULTS_4_2(79)<=signed(MULTS_3_2(79)(PERCISION) & MULTS_3_2(79)(PERCISION downto 1))+signed(MULTS_3_3(79)(PERCISION) & MULTS_3_3(79)(PERCISION downto 1));
			MULTS_4_2(80)<=signed(MULTS_3_2(80)(PERCISION) & MULTS_3_2(80)(PERCISION downto 1))+signed(MULTS_3_3(80)(PERCISION) & MULTS_3_3(80)(PERCISION downto 1));
			MULTS_4_2(81)<=signed(MULTS_3_2(81)(PERCISION) & MULTS_3_2(81)(PERCISION downto 1))+signed(MULTS_3_3(81)(PERCISION) & MULTS_3_3(81)(PERCISION downto 1));
			MULTS_4_2(82)<=signed(MULTS_3_2(82)(PERCISION) & MULTS_3_2(82)(PERCISION downto 1))+signed(MULTS_3_3(82)(PERCISION) & MULTS_3_3(82)(PERCISION downto 1));
			MULTS_4_2(83)<=signed(MULTS_3_2(83)(PERCISION) & MULTS_3_2(83)(PERCISION downto 1))+signed(MULTS_3_3(83)(PERCISION) & MULTS_3_3(83)(PERCISION downto 1));

			MULTS_4_3(0)<=signed(MULTS_3_4(0)(PERCISION) & MULTS_3_4(0)(PERCISION downto 1))+signed(MULTS_3_5(0)(PERCISION) & MULTS_3_5(0)(PERCISION downto 1));
			MULTS_4_3(1)<=signed(MULTS_3_4(1)(PERCISION) & MULTS_3_4(1)(PERCISION downto 1))+signed(MULTS_3_5(1)(PERCISION) & MULTS_3_5(1)(PERCISION downto 1));
			MULTS_4_3(2)<=signed(MULTS_3_4(2)(PERCISION) & MULTS_3_4(2)(PERCISION downto 1))+signed(MULTS_3_5(2)(PERCISION) & MULTS_3_5(2)(PERCISION downto 1));
			MULTS_4_3(3)<=signed(MULTS_3_4(3)(PERCISION) & MULTS_3_4(3)(PERCISION downto 1))+signed(MULTS_3_5(3)(PERCISION) & MULTS_3_5(3)(PERCISION downto 1));
			MULTS_4_3(4)<=signed(MULTS_3_4(4)(PERCISION) & MULTS_3_4(4)(PERCISION downto 1))+signed(MULTS_3_5(4)(PERCISION) & MULTS_3_5(4)(PERCISION downto 1));
			MULTS_4_3(5)<=signed(MULTS_3_4(5)(PERCISION) & MULTS_3_4(5)(PERCISION downto 1))+signed(MULTS_3_5(5)(PERCISION) & MULTS_3_5(5)(PERCISION downto 1));
			MULTS_4_3(6)<=signed(MULTS_3_4(6)(PERCISION) & MULTS_3_4(6)(PERCISION downto 1))+signed(MULTS_3_5(6)(PERCISION) & MULTS_3_5(6)(PERCISION downto 1));
			MULTS_4_3(7)<=signed(MULTS_3_4(7)(PERCISION) & MULTS_3_4(7)(PERCISION downto 1))+signed(MULTS_3_5(7)(PERCISION) & MULTS_3_5(7)(PERCISION downto 1));
			MULTS_4_3(8)<=signed(MULTS_3_4(8)(PERCISION) & MULTS_3_4(8)(PERCISION downto 1))+signed(MULTS_3_5(8)(PERCISION) & MULTS_3_5(8)(PERCISION downto 1));
			MULTS_4_3(9)<=signed(MULTS_3_4(9)(PERCISION) & MULTS_3_4(9)(PERCISION downto 1))+signed(MULTS_3_5(9)(PERCISION) & MULTS_3_5(9)(PERCISION downto 1));
			MULTS_4_3(10)<=signed(MULTS_3_4(10)(PERCISION) & MULTS_3_4(10)(PERCISION downto 1))+signed(MULTS_3_5(10)(PERCISION) & MULTS_3_5(10)(PERCISION downto 1));
			MULTS_4_3(11)<=signed(MULTS_3_4(11)(PERCISION) & MULTS_3_4(11)(PERCISION downto 1))+signed(MULTS_3_5(11)(PERCISION) & MULTS_3_5(11)(PERCISION downto 1));
			MULTS_4_3(12)<=signed(MULTS_3_4(12)(PERCISION) & MULTS_3_4(12)(PERCISION downto 1))+signed(MULTS_3_5(12)(PERCISION) & MULTS_3_5(12)(PERCISION downto 1));
			MULTS_4_3(13)<=signed(MULTS_3_4(13)(PERCISION) & MULTS_3_4(13)(PERCISION downto 1))+signed(MULTS_3_5(13)(PERCISION) & MULTS_3_5(13)(PERCISION downto 1));
			MULTS_4_3(14)<=signed(MULTS_3_4(14)(PERCISION) & MULTS_3_4(14)(PERCISION downto 1))+signed(MULTS_3_5(14)(PERCISION) & MULTS_3_5(14)(PERCISION downto 1));
			MULTS_4_3(15)<=signed(MULTS_3_4(15)(PERCISION) & MULTS_3_4(15)(PERCISION downto 1))+signed(MULTS_3_5(15)(PERCISION) & MULTS_3_5(15)(PERCISION downto 1));
			MULTS_4_3(16)<=signed(MULTS_3_4(16)(PERCISION) & MULTS_3_4(16)(PERCISION downto 1))+signed(MULTS_3_5(16)(PERCISION) & MULTS_3_5(16)(PERCISION downto 1));
			MULTS_4_3(17)<=signed(MULTS_3_4(17)(PERCISION) & MULTS_3_4(17)(PERCISION downto 1))+signed(MULTS_3_5(17)(PERCISION) & MULTS_3_5(17)(PERCISION downto 1));
			MULTS_4_3(18)<=signed(MULTS_3_4(18)(PERCISION) & MULTS_3_4(18)(PERCISION downto 1))+signed(MULTS_3_5(18)(PERCISION) & MULTS_3_5(18)(PERCISION downto 1));
			MULTS_4_3(19)<=signed(MULTS_3_4(19)(PERCISION) & MULTS_3_4(19)(PERCISION downto 1))+signed(MULTS_3_5(19)(PERCISION) & MULTS_3_5(19)(PERCISION downto 1));
			MULTS_4_3(20)<=signed(MULTS_3_4(20)(PERCISION) & MULTS_3_4(20)(PERCISION downto 1))+signed(MULTS_3_5(20)(PERCISION) & MULTS_3_5(20)(PERCISION downto 1));
			MULTS_4_3(21)<=signed(MULTS_3_4(21)(PERCISION) & MULTS_3_4(21)(PERCISION downto 1))+signed(MULTS_3_5(21)(PERCISION) & MULTS_3_5(21)(PERCISION downto 1));
			MULTS_4_3(22)<=signed(MULTS_3_4(22)(PERCISION) & MULTS_3_4(22)(PERCISION downto 1))+signed(MULTS_3_5(22)(PERCISION) & MULTS_3_5(22)(PERCISION downto 1));
			MULTS_4_3(23)<=signed(MULTS_3_4(23)(PERCISION) & MULTS_3_4(23)(PERCISION downto 1))+signed(MULTS_3_5(23)(PERCISION) & MULTS_3_5(23)(PERCISION downto 1));
			MULTS_4_3(24)<=signed(MULTS_3_4(24)(PERCISION) & MULTS_3_4(24)(PERCISION downto 1))+signed(MULTS_3_5(24)(PERCISION) & MULTS_3_5(24)(PERCISION downto 1));
			MULTS_4_3(25)<=signed(MULTS_3_4(25)(PERCISION) & MULTS_3_4(25)(PERCISION downto 1))+signed(MULTS_3_5(25)(PERCISION) & MULTS_3_5(25)(PERCISION downto 1));
			MULTS_4_3(26)<=signed(MULTS_3_4(26)(PERCISION) & MULTS_3_4(26)(PERCISION downto 1))+signed(MULTS_3_5(26)(PERCISION) & MULTS_3_5(26)(PERCISION downto 1));
			MULTS_4_3(27)<=signed(MULTS_3_4(27)(PERCISION) & MULTS_3_4(27)(PERCISION downto 1))+signed(MULTS_3_5(27)(PERCISION) & MULTS_3_5(27)(PERCISION downto 1));
			MULTS_4_3(28)<=signed(MULTS_3_4(28)(PERCISION) & MULTS_3_4(28)(PERCISION downto 1))+signed(MULTS_3_5(28)(PERCISION) & MULTS_3_5(28)(PERCISION downto 1));
			MULTS_4_3(29)<=signed(MULTS_3_4(29)(PERCISION) & MULTS_3_4(29)(PERCISION downto 1))+signed(MULTS_3_5(29)(PERCISION) & MULTS_3_5(29)(PERCISION downto 1));
			MULTS_4_3(30)<=signed(MULTS_3_4(30)(PERCISION) & MULTS_3_4(30)(PERCISION downto 1))+signed(MULTS_3_5(30)(PERCISION) & MULTS_3_5(30)(PERCISION downto 1));
			MULTS_4_3(31)<=signed(MULTS_3_4(31)(PERCISION) & MULTS_3_4(31)(PERCISION downto 1))+signed(MULTS_3_5(31)(PERCISION) & MULTS_3_5(31)(PERCISION downto 1));
			MULTS_4_3(32)<=signed(MULTS_3_4(32)(PERCISION) & MULTS_3_4(32)(PERCISION downto 1))+signed(MULTS_3_5(32)(PERCISION) & MULTS_3_5(32)(PERCISION downto 1));
			MULTS_4_3(33)<=signed(MULTS_3_4(33)(PERCISION) & MULTS_3_4(33)(PERCISION downto 1))+signed(MULTS_3_5(33)(PERCISION) & MULTS_3_5(33)(PERCISION downto 1));
			MULTS_4_3(34)<=signed(MULTS_3_4(34)(PERCISION) & MULTS_3_4(34)(PERCISION downto 1))+signed(MULTS_3_5(34)(PERCISION) & MULTS_3_5(34)(PERCISION downto 1));
			MULTS_4_3(35)<=signed(MULTS_3_4(35)(PERCISION) & MULTS_3_4(35)(PERCISION downto 1))+signed(MULTS_3_5(35)(PERCISION) & MULTS_3_5(35)(PERCISION downto 1));
			MULTS_4_3(36)<=signed(MULTS_3_4(36)(PERCISION) & MULTS_3_4(36)(PERCISION downto 1))+signed(MULTS_3_5(36)(PERCISION) & MULTS_3_5(36)(PERCISION downto 1));
			MULTS_4_3(37)<=signed(MULTS_3_4(37)(PERCISION) & MULTS_3_4(37)(PERCISION downto 1))+signed(MULTS_3_5(37)(PERCISION) & MULTS_3_5(37)(PERCISION downto 1));
			MULTS_4_3(38)<=signed(MULTS_3_4(38)(PERCISION) & MULTS_3_4(38)(PERCISION downto 1))+signed(MULTS_3_5(38)(PERCISION) & MULTS_3_5(38)(PERCISION downto 1));
			MULTS_4_3(39)<=signed(MULTS_3_4(39)(PERCISION) & MULTS_3_4(39)(PERCISION downto 1))+signed(MULTS_3_5(39)(PERCISION) & MULTS_3_5(39)(PERCISION downto 1));
			MULTS_4_3(40)<=signed(MULTS_3_4(40)(PERCISION) & MULTS_3_4(40)(PERCISION downto 1))+signed(MULTS_3_5(40)(PERCISION) & MULTS_3_5(40)(PERCISION downto 1));
			MULTS_4_3(41)<=signed(MULTS_3_4(41)(PERCISION) & MULTS_3_4(41)(PERCISION downto 1))+signed(MULTS_3_5(41)(PERCISION) & MULTS_3_5(41)(PERCISION downto 1));
			MULTS_4_3(42)<=signed(MULTS_3_4(42)(PERCISION) & MULTS_3_4(42)(PERCISION downto 1))+signed(MULTS_3_5(42)(PERCISION) & MULTS_3_5(42)(PERCISION downto 1));
			MULTS_4_3(43)<=signed(MULTS_3_4(43)(PERCISION) & MULTS_3_4(43)(PERCISION downto 1))+signed(MULTS_3_5(43)(PERCISION) & MULTS_3_5(43)(PERCISION downto 1));
			MULTS_4_3(44)<=signed(MULTS_3_4(44)(PERCISION) & MULTS_3_4(44)(PERCISION downto 1))+signed(MULTS_3_5(44)(PERCISION) & MULTS_3_5(44)(PERCISION downto 1));
			MULTS_4_3(45)<=signed(MULTS_3_4(45)(PERCISION) & MULTS_3_4(45)(PERCISION downto 1))+signed(MULTS_3_5(45)(PERCISION) & MULTS_3_5(45)(PERCISION downto 1));
			MULTS_4_3(46)<=signed(MULTS_3_4(46)(PERCISION) & MULTS_3_4(46)(PERCISION downto 1))+signed(MULTS_3_5(46)(PERCISION) & MULTS_3_5(46)(PERCISION downto 1));
			MULTS_4_3(47)<=signed(MULTS_3_4(47)(PERCISION) & MULTS_3_4(47)(PERCISION downto 1))+signed(MULTS_3_5(47)(PERCISION) & MULTS_3_5(47)(PERCISION downto 1));
			MULTS_4_3(48)<=signed(MULTS_3_4(48)(PERCISION) & MULTS_3_4(48)(PERCISION downto 1))+signed(MULTS_3_5(48)(PERCISION) & MULTS_3_5(48)(PERCISION downto 1));
			MULTS_4_3(49)<=signed(MULTS_3_4(49)(PERCISION) & MULTS_3_4(49)(PERCISION downto 1))+signed(MULTS_3_5(49)(PERCISION) & MULTS_3_5(49)(PERCISION downto 1));
			MULTS_4_3(50)<=signed(MULTS_3_4(50)(PERCISION) & MULTS_3_4(50)(PERCISION downto 1))+signed(MULTS_3_5(50)(PERCISION) & MULTS_3_5(50)(PERCISION downto 1));
			MULTS_4_3(51)<=signed(MULTS_3_4(51)(PERCISION) & MULTS_3_4(51)(PERCISION downto 1))+signed(MULTS_3_5(51)(PERCISION) & MULTS_3_5(51)(PERCISION downto 1));
			MULTS_4_3(52)<=signed(MULTS_3_4(52)(PERCISION) & MULTS_3_4(52)(PERCISION downto 1))+signed(MULTS_3_5(52)(PERCISION) & MULTS_3_5(52)(PERCISION downto 1));
			MULTS_4_3(53)<=signed(MULTS_3_4(53)(PERCISION) & MULTS_3_4(53)(PERCISION downto 1))+signed(MULTS_3_5(53)(PERCISION) & MULTS_3_5(53)(PERCISION downto 1));
			MULTS_4_3(54)<=signed(MULTS_3_4(54)(PERCISION) & MULTS_3_4(54)(PERCISION downto 1))+signed(MULTS_3_5(54)(PERCISION) & MULTS_3_5(54)(PERCISION downto 1));
			MULTS_4_3(55)<=signed(MULTS_3_4(55)(PERCISION) & MULTS_3_4(55)(PERCISION downto 1))+signed(MULTS_3_5(55)(PERCISION) & MULTS_3_5(55)(PERCISION downto 1));
			MULTS_4_3(56)<=signed(MULTS_3_4(56)(PERCISION) & MULTS_3_4(56)(PERCISION downto 1))+signed(MULTS_3_5(56)(PERCISION) & MULTS_3_5(56)(PERCISION downto 1));
			MULTS_4_3(57)<=signed(MULTS_3_4(57)(PERCISION) & MULTS_3_4(57)(PERCISION downto 1))+signed(MULTS_3_5(57)(PERCISION) & MULTS_3_5(57)(PERCISION downto 1));
			MULTS_4_3(58)<=signed(MULTS_3_4(58)(PERCISION) & MULTS_3_4(58)(PERCISION downto 1))+signed(MULTS_3_5(58)(PERCISION) & MULTS_3_5(58)(PERCISION downto 1));
			MULTS_4_3(59)<=signed(MULTS_3_4(59)(PERCISION) & MULTS_3_4(59)(PERCISION downto 1))+signed(MULTS_3_5(59)(PERCISION) & MULTS_3_5(59)(PERCISION downto 1));
			MULTS_4_3(60)<=signed(MULTS_3_4(60)(PERCISION) & MULTS_3_4(60)(PERCISION downto 1))+signed(MULTS_3_5(60)(PERCISION) & MULTS_3_5(60)(PERCISION downto 1));
			MULTS_4_3(61)<=signed(MULTS_3_4(61)(PERCISION) & MULTS_3_4(61)(PERCISION downto 1))+signed(MULTS_3_5(61)(PERCISION) & MULTS_3_5(61)(PERCISION downto 1));
			MULTS_4_3(62)<=signed(MULTS_3_4(62)(PERCISION) & MULTS_3_4(62)(PERCISION downto 1))+signed(MULTS_3_5(62)(PERCISION) & MULTS_3_5(62)(PERCISION downto 1));
			MULTS_4_3(63)<=signed(MULTS_3_4(63)(PERCISION) & MULTS_3_4(63)(PERCISION downto 1))+signed(MULTS_3_5(63)(PERCISION) & MULTS_3_5(63)(PERCISION downto 1));
			MULTS_4_3(64)<=signed(MULTS_3_4(64)(PERCISION) & MULTS_3_4(64)(PERCISION downto 1))+signed(MULTS_3_5(64)(PERCISION) & MULTS_3_5(64)(PERCISION downto 1));
			MULTS_4_3(65)<=signed(MULTS_3_4(65)(PERCISION) & MULTS_3_4(65)(PERCISION downto 1))+signed(MULTS_3_5(65)(PERCISION) & MULTS_3_5(65)(PERCISION downto 1));
			MULTS_4_3(66)<=signed(MULTS_3_4(66)(PERCISION) & MULTS_3_4(66)(PERCISION downto 1))+signed(MULTS_3_5(66)(PERCISION) & MULTS_3_5(66)(PERCISION downto 1));
			MULTS_4_3(67)<=signed(MULTS_3_4(67)(PERCISION) & MULTS_3_4(67)(PERCISION downto 1))+signed(MULTS_3_5(67)(PERCISION) & MULTS_3_5(67)(PERCISION downto 1));
			MULTS_4_3(68)<=signed(MULTS_3_4(68)(PERCISION) & MULTS_3_4(68)(PERCISION downto 1))+signed(MULTS_3_5(68)(PERCISION) & MULTS_3_5(68)(PERCISION downto 1));
			MULTS_4_3(69)<=signed(MULTS_3_4(69)(PERCISION) & MULTS_3_4(69)(PERCISION downto 1))+signed(MULTS_3_5(69)(PERCISION) & MULTS_3_5(69)(PERCISION downto 1));
			MULTS_4_3(70)<=signed(MULTS_3_4(70)(PERCISION) & MULTS_3_4(70)(PERCISION downto 1))+signed(MULTS_3_5(70)(PERCISION) & MULTS_3_5(70)(PERCISION downto 1));
			MULTS_4_3(71)<=signed(MULTS_3_4(71)(PERCISION) & MULTS_3_4(71)(PERCISION downto 1))+signed(MULTS_3_5(71)(PERCISION) & MULTS_3_5(71)(PERCISION downto 1));
			MULTS_4_3(72)<=signed(MULTS_3_4(72)(PERCISION) & MULTS_3_4(72)(PERCISION downto 1))+signed(MULTS_3_5(72)(PERCISION) & MULTS_3_5(72)(PERCISION downto 1));
			MULTS_4_3(73)<=signed(MULTS_3_4(73)(PERCISION) & MULTS_3_4(73)(PERCISION downto 1))+signed(MULTS_3_5(73)(PERCISION) & MULTS_3_5(73)(PERCISION downto 1));
			MULTS_4_3(74)<=signed(MULTS_3_4(74)(PERCISION) & MULTS_3_4(74)(PERCISION downto 1))+signed(MULTS_3_5(74)(PERCISION) & MULTS_3_5(74)(PERCISION downto 1));
			MULTS_4_3(75)<=signed(MULTS_3_4(75)(PERCISION) & MULTS_3_4(75)(PERCISION downto 1))+signed(MULTS_3_5(75)(PERCISION) & MULTS_3_5(75)(PERCISION downto 1));
			MULTS_4_3(76)<=signed(MULTS_3_4(76)(PERCISION) & MULTS_3_4(76)(PERCISION downto 1))+signed(MULTS_3_5(76)(PERCISION) & MULTS_3_5(76)(PERCISION downto 1));
			MULTS_4_3(77)<=signed(MULTS_3_4(77)(PERCISION) & MULTS_3_4(77)(PERCISION downto 1))+signed(MULTS_3_5(77)(PERCISION) & MULTS_3_5(77)(PERCISION downto 1));
			MULTS_4_3(78)<=signed(MULTS_3_4(78)(PERCISION) & MULTS_3_4(78)(PERCISION downto 1))+signed(MULTS_3_5(78)(PERCISION) & MULTS_3_5(78)(PERCISION downto 1));
			MULTS_4_3(79)<=signed(MULTS_3_4(79)(PERCISION) & MULTS_3_4(79)(PERCISION downto 1))+signed(MULTS_3_5(79)(PERCISION) & MULTS_3_5(79)(PERCISION downto 1));
			MULTS_4_3(80)<=signed(MULTS_3_4(80)(PERCISION) & MULTS_3_4(80)(PERCISION downto 1))+signed(MULTS_3_5(80)(PERCISION) & MULTS_3_5(80)(PERCISION downto 1));
			MULTS_4_3(81)<=signed(MULTS_3_4(81)(PERCISION) & MULTS_3_4(81)(PERCISION downto 1))+signed(MULTS_3_5(81)(PERCISION) & MULTS_3_5(81)(PERCISION downto 1));
			MULTS_4_3(82)<=signed(MULTS_3_4(82)(PERCISION) & MULTS_3_4(82)(PERCISION downto 1))+signed(MULTS_3_5(82)(PERCISION) & MULTS_3_5(82)(PERCISION downto 1));
			MULTS_4_3(83)<=signed(MULTS_3_4(83)(PERCISION) & MULTS_3_4(83)(PERCISION downto 1))+signed(MULTS_3_5(83)(PERCISION) & MULTS_3_5(83)(PERCISION downto 1));

			MULTS_4_4(0)<=signed(MULTS_3_6(0)(PERCISION) & MULTS_3_6(0)(PERCISION downto 1))+signed(MULTS_3_7(0)(PERCISION) & MULTS_3_7(0)(PERCISION downto 1));
			MULTS_4_4(1)<=signed(MULTS_3_6(1)(PERCISION) & MULTS_3_6(1)(PERCISION downto 1))+signed(MULTS_3_7(1)(PERCISION) & MULTS_3_7(1)(PERCISION downto 1));
			MULTS_4_4(2)<=signed(MULTS_3_6(2)(PERCISION) & MULTS_3_6(2)(PERCISION downto 1))+signed(MULTS_3_7(2)(PERCISION) & MULTS_3_7(2)(PERCISION downto 1));
			MULTS_4_4(3)<=signed(MULTS_3_6(3)(PERCISION) & MULTS_3_6(3)(PERCISION downto 1))+signed(MULTS_3_7(3)(PERCISION) & MULTS_3_7(3)(PERCISION downto 1));
			MULTS_4_4(4)<=signed(MULTS_3_6(4)(PERCISION) & MULTS_3_6(4)(PERCISION downto 1))+signed(MULTS_3_7(4)(PERCISION) & MULTS_3_7(4)(PERCISION downto 1));
			MULTS_4_4(5)<=signed(MULTS_3_6(5)(PERCISION) & MULTS_3_6(5)(PERCISION downto 1))+signed(MULTS_3_7(5)(PERCISION) & MULTS_3_7(5)(PERCISION downto 1));
			MULTS_4_4(6)<=signed(MULTS_3_6(6)(PERCISION) & MULTS_3_6(6)(PERCISION downto 1))+signed(MULTS_3_7(6)(PERCISION) & MULTS_3_7(6)(PERCISION downto 1));
			MULTS_4_4(7)<=signed(MULTS_3_6(7)(PERCISION) & MULTS_3_6(7)(PERCISION downto 1))+signed(MULTS_3_7(7)(PERCISION) & MULTS_3_7(7)(PERCISION downto 1));
			MULTS_4_4(8)<=signed(MULTS_3_6(8)(PERCISION) & MULTS_3_6(8)(PERCISION downto 1))+signed(MULTS_3_7(8)(PERCISION) & MULTS_3_7(8)(PERCISION downto 1));
			MULTS_4_4(9)<=signed(MULTS_3_6(9)(PERCISION) & MULTS_3_6(9)(PERCISION downto 1))+signed(MULTS_3_7(9)(PERCISION) & MULTS_3_7(9)(PERCISION downto 1));
			MULTS_4_4(10)<=signed(MULTS_3_6(10)(PERCISION) & MULTS_3_6(10)(PERCISION downto 1))+signed(MULTS_3_7(10)(PERCISION) & MULTS_3_7(10)(PERCISION downto 1));
			MULTS_4_4(11)<=signed(MULTS_3_6(11)(PERCISION) & MULTS_3_6(11)(PERCISION downto 1))+signed(MULTS_3_7(11)(PERCISION) & MULTS_3_7(11)(PERCISION downto 1));
			MULTS_4_4(12)<=signed(MULTS_3_6(12)(PERCISION) & MULTS_3_6(12)(PERCISION downto 1))+signed(MULTS_3_7(12)(PERCISION) & MULTS_3_7(12)(PERCISION downto 1));
			MULTS_4_4(13)<=signed(MULTS_3_6(13)(PERCISION) & MULTS_3_6(13)(PERCISION downto 1))+signed(MULTS_3_7(13)(PERCISION) & MULTS_3_7(13)(PERCISION downto 1));
			MULTS_4_4(14)<=signed(MULTS_3_6(14)(PERCISION) & MULTS_3_6(14)(PERCISION downto 1))+signed(MULTS_3_7(14)(PERCISION) & MULTS_3_7(14)(PERCISION downto 1));
			MULTS_4_4(15)<=signed(MULTS_3_6(15)(PERCISION) & MULTS_3_6(15)(PERCISION downto 1))+signed(MULTS_3_7(15)(PERCISION) & MULTS_3_7(15)(PERCISION downto 1));
			MULTS_4_4(16)<=signed(MULTS_3_6(16)(PERCISION) & MULTS_3_6(16)(PERCISION downto 1))+signed(MULTS_3_7(16)(PERCISION) & MULTS_3_7(16)(PERCISION downto 1));
			MULTS_4_4(17)<=signed(MULTS_3_6(17)(PERCISION) & MULTS_3_6(17)(PERCISION downto 1))+signed(MULTS_3_7(17)(PERCISION) & MULTS_3_7(17)(PERCISION downto 1));
			MULTS_4_4(18)<=signed(MULTS_3_6(18)(PERCISION) & MULTS_3_6(18)(PERCISION downto 1))+signed(MULTS_3_7(18)(PERCISION) & MULTS_3_7(18)(PERCISION downto 1));
			MULTS_4_4(19)<=signed(MULTS_3_6(19)(PERCISION) & MULTS_3_6(19)(PERCISION downto 1))+signed(MULTS_3_7(19)(PERCISION) & MULTS_3_7(19)(PERCISION downto 1));
			MULTS_4_4(20)<=signed(MULTS_3_6(20)(PERCISION) & MULTS_3_6(20)(PERCISION downto 1))+signed(MULTS_3_7(20)(PERCISION) & MULTS_3_7(20)(PERCISION downto 1));
			MULTS_4_4(21)<=signed(MULTS_3_6(21)(PERCISION) & MULTS_3_6(21)(PERCISION downto 1))+signed(MULTS_3_7(21)(PERCISION) & MULTS_3_7(21)(PERCISION downto 1));
			MULTS_4_4(22)<=signed(MULTS_3_6(22)(PERCISION) & MULTS_3_6(22)(PERCISION downto 1))+signed(MULTS_3_7(22)(PERCISION) & MULTS_3_7(22)(PERCISION downto 1));
			MULTS_4_4(23)<=signed(MULTS_3_6(23)(PERCISION) & MULTS_3_6(23)(PERCISION downto 1))+signed(MULTS_3_7(23)(PERCISION) & MULTS_3_7(23)(PERCISION downto 1));
			MULTS_4_4(24)<=signed(MULTS_3_6(24)(PERCISION) & MULTS_3_6(24)(PERCISION downto 1))+signed(MULTS_3_7(24)(PERCISION) & MULTS_3_7(24)(PERCISION downto 1));
			MULTS_4_4(25)<=signed(MULTS_3_6(25)(PERCISION) & MULTS_3_6(25)(PERCISION downto 1))+signed(MULTS_3_7(25)(PERCISION) & MULTS_3_7(25)(PERCISION downto 1));
			MULTS_4_4(26)<=signed(MULTS_3_6(26)(PERCISION) & MULTS_3_6(26)(PERCISION downto 1))+signed(MULTS_3_7(26)(PERCISION) & MULTS_3_7(26)(PERCISION downto 1));
			MULTS_4_4(27)<=signed(MULTS_3_6(27)(PERCISION) & MULTS_3_6(27)(PERCISION downto 1))+signed(MULTS_3_7(27)(PERCISION) & MULTS_3_7(27)(PERCISION downto 1));
			MULTS_4_4(28)<=signed(MULTS_3_6(28)(PERCISION) & MULTS_3_6(28)(PERCISION downto 1))+signed(MULTS_3_7(28)(PERCISION) & MULTS_3_7(28)(PERCISION downto 1));
			MULTS_4_4(29)<=signed(MULTS_3_6(29)(PERCISION) & MULTS_3_6(29)(PERCISION downto 1))+signed(MULTS_3_7(29)(PERCISION) & MULTS_3_7(29)(PERCISION downto 1));
			MULTS_4_4(30)<=signed(MULTS_3_6(30)(PERCISION) & MULTS_3_6(30)(PERCISION downto 1))+signed(MULTS_3_7(30)(PERCISION) & MULTS_3_7(30)(PERCISION downto 1));
			MULTS_4_4(31)<=signed(MULTS_3_6(31)(PERCISION) & MULTS_3_6(31)(PERCISION downto 1))+signed(MULTS_3_7(31)(PERCISION) & MULTS_3_7(31)(PERCISION downto 1));
			MULTS_4_4(32)<=signed(MULTS_3_6(32)(PERCISION) & MULTS_3_6(32)(PERCISION downto 1))+signed(MULTS_3_7(32)(PERCISION) & MULTS_3_7(32)(PERCISION downto 1));
			MULTS_4_4(33)<=signed(MULTS_3_6(33)(PERCISION) & MULTS_3_6(33)(PERCISION downto 1))+signed(MULTS_3_7(33)(PERCISION) & MULTS_3_7(33)(PERCISION downto 1));
			MULTS_4_4(34)<=signed(MULTS_3_6(34)(PERCISION) & MULTS_3_6(34)(PERCISION downto 1))+signed(MULTS_3_7(34)(PERCISION) & MULTS_3_7(34)(PERCISION downto 1));
			MULTS_4_4(35)<=signed(MULTS_3_6(35)(PERCISION) & MULTS_3_6(35)(PERCISION downto 1))+signed(MULTS_3_7(35)(PERCISION) & MULTS_3_7(35)(PERCISION downto 1));
			MULTS_4_4(36)<=signed(MULTS_3_6(36)(PERCISION) & MULTS_3_6(36)(PERCISION downto 1))+signed(MULTS_3_7(36)(PERCISION) & MULTS_3_7(36)(PERCISION downto 1));
			MULTS_4_4(37)<=signed(MULTS_3_6(37)(PERCISION) & MULTS_3_6(37)(PERCISION downto 1))+signed(MULTS_3_7(37)(PERCISION) & MULTS_3_7(37)(PERCISION downto 1));
			MULTS_4_4(38)<=signed(MULTS_3_6(38)(PERCISION) & MULTS_3_6(38)(PERCISION downto 1))+signed(MULTS_3_7(38)(PERCISION) & MULTS_3_7(38)(PERCISION downto 1));
			MULTS_4_4(39)<=signed(MULTS_3_6(39)(PERCISION) & MULTS_3_6(39)(PERCISION downto 1))+signed(MULTS_3_7(39)(PERCISION) & MULTS_3_7(39)(PERCISION downto 1));
			MULTS_4_4(40)<=signed(MULTS_3_6(40)(PERCISION) & MULTS_3_6(40)(PERCISION downto 1))+signed(MULTS_3_7(40)(PERCISION) & MULTS_3_7(40)(PERCISION downto 1));
			MULTS_4_4(41)<=signed(MULTS_3_6(41)(PERCISION) & MULTS_3_6(41)(PERCISION downto 1))+signed(MULTS_3_7(41)(PERCISION) & MULTS_3_7(41)(PERCISION downto 1));
			MULTS_4_4(42)<=signed(MULTS_3_6(42)(PERCISION) & MULTS_3_6(42)(PERCISION downto 1))+signed(MULTS_3_7(42)(PERCISION) & MULTS_3_7(42)(PERCISION downto 1));
			MULTS_4_4(43)<=signed(MULTS_3_6(43)(PERCISION) & MULTS_3_6(43)(PERCISION downto 1))+signed(MULTS_3_7(43)(PERCISION) & MULTS_3_7(43)(PERCISION downto 1));
			MULTS_4_4(44)<=signed(MULTS_3_6(44)(PERCISION) & MULTS_3_6(44)(PERCISION downto 1))+signed(MULTS_3_7(44)(PERCISION) & MULTS_3_7(44)(PERCISION downto 1));
			MULTS_4_4(45)<=signed(MULTS_3_6(45)(PERCISION) & MULTS_3_6(45)(PERCISION downto 1))+signed(MULTS_3_7(45)(PERCISION) & MULTS_3_7(45)(PERCISION downto 1));
			MULTS_4_4(46)<=signed(MULTS_3_6(46)(PERCISION) & MULTS_3_6(46)(PERCISION downto 1))+signed(MULTS_3_7(46)(PERCISION) & MULTS_3_7(46)(PERCISION downto 1));
			MULTS_4_4(47)<=signed(MULTS_3_6(47)(PERCISION) & MULTS_3_6(47)(PERCISION downto 1))+signed(MULTS_3_7(47)(PERCISION) & MULTS_3_7(47)(PERCISION downto 1));
			MULTS_4_4(48)<=signed(MULTS_3_6(48)(PERCISION) & MULTS_3_6(48)(PERCISION downto 1))+signed(MULTS_3_7(48)(PERCISION) & MULTS_3_7(48)(PERCISION downto 1));
			MULTS_4_4(49)<=signed(MULTS_3_6(49)(PERCISION) & MULTS_3_6(49)(PERCISION downto 1))+signed(MULTS_3_7(49)(PERCISION) & MULTS_3_7(49)(PERCISION downto 1));
			MULTS_4_4(50)<=signed(MULTS_3_6(50)(PERCISION) & MULTS_3_6(50)(PERCISION downto 1))+signed(MULTS_3_7(50)(PERCISION) & MULTS_3_7(50)(PERCISION downto 1));
			MULTS_4_4(51)<=signed(MULTS_3_6(51)(PERCISION) & MULTS_3_6(51)(PERCISION downto 1))+signed(MULTS_3_7(51)(PERCISION) & MULTS_3_7(51)(PERCISION downto 1));
			MULTS_4_4(52)<=signed(MULTS_3_6(52)(PERCISION) & MULTS_3_6(52)(PERCISION downto 1))+signed(MULTS_3_7(52)(PERCISION) & MULTS_3_7(52)(PERCISION downto 1));
			MULTS_4_4(53)<=signed(MULTS_3_6(53)(PERCISION) & MULTS_3_6(53)(PERCISION downto 1))+signed(MULTS_3_7(53)(PERCISION) & MULTS_3_7(53)(PERCISION downto 1));
			MULTS_4_4(54)<=signed(MULTS_3_6(54)(PERCISION) & MULTS_3_6(54)(PERCISION downto 1))+signed(MULTS_3_7(54)(PERCISION) & MULTS_3_7(54)(PERCISION downto 1));
			MULTS_4_4(55)<=signed(MULTS_3_6(55)(PERCISION) & MULTS_3_6(55)(PERCISION downto 1))+signed(MULTS_3_7(55)(PERCISION) & MULTS_3_7(55)(PERCISION downto 1));
			MULTS_4_4(56)<=signed(MULTS_3_6(56)(PERCISION) & MULTS_3_6(56)(PERCISION downto 1))+signed(MULTS_3_7(56)(PERCISION) & MULTS_3_7(56)(PERCISION downto 1));
			MULTS_4_4(57)<=signed(MULTS_3_6(57)(PERCISION) & MULTS_3_6(57)(PERCISION downto 1))+signed(MULTS_3_7(57)(PERCISION) & MULTS_3_7(57)(PERCISION downto 1));
			MULTS_4_4(58)<=signed(MULTS_3_6(58)(PERCISION) & MULTS_3_6(58)(PERCISION downto 1))+signed(MULTS_3_7(58)(PERCISION) & MULTS_3_7(58)(PERCISION downto 1));
			MULTS_4_4(59)<=signed(MULTS_3_6(59)(PERCISION) & MULTS_3_6(59)(PERCISION downto 1))+signed(MULTS_3_7(59)(PERCISION) & MULTS_3_7(59)(PERCISION downto 1));
			MULTS_4_4(60)<=signed(MULTS_3_6(60)(PERCISION) & MULTS_3_6(60)(PERCISION downto 1))+signed(MULTS_3_7(60)(PERCISION) & MULTS_3_7(60)(PERCISION downto 1));
			MULTS_4_4(61)<=signed(MULTS_3_6(61)(PERCISION) & MULTS_3_6(61)(PERCISION downto 1))+signed(MULTS_3_7(61)(PERCISION) & MULTS_3_7(61)(PERCISION downto 1));
			MULTS_4_4(62)<=signed(MULTS_3_6(62)(PERCISION) & MULTS_3_6(62)(PERCISION downto 1))+signed(MULTS_3_7(62)(PERCISION) & MULTS_3_7(62)(PERCISION downto 1));
			MULTS_4_4(63)<=signed(MULTS_3_6(63)(PERCISION) & MULTS_3_6(63)(PERCISION downto 1))+signed(MULTS_3_7(63)(PERCISION) & MULTS_3_7(63)(PERCISION downto 1));
			MULTS_4_4(64)<=signed(MULTS_3_6(64)(PERCISION) & MULTS_3_6(64)(PERCISION downto 1))+signed(MULTS_3_7(64)(PERCISION) & MULTS_3_7(64)(PERCISION downto 1));
			MULTS_4_4(65)<=signed(MULTS_3_6(65)(PERCISION) & MULTS_3_6(65)(PERCISION downto 1))+signed(MULTS_3_7(65)(PERCISION) & MULTS_3_7(65)(PERCISION downto 1));
			MULTS_4_4(66)<=signed(MULTS_3_6(66)(PERCISION) & MULTS_3_6(66)(PERCISION downto 1))+signed(MULTS_3_7(66)(PERCISION) & MULTS_3_7(66)(PERCISION downto 1));
			MULTS_4_4(67)<=signed(MULTS_3_6(67)(PERCISION) & MULTS_3_6(67)(PERCISION downto 1))+signed(MULTS_3_7(67)(PERCISION) & MULTS_3_7(67)(PERCISION downto 1));
			MULTS_4_4(68)<=signed(MULTS_3_6(68)(PERCISION) & MULTS_3_6(68)(PERCISION downto 1))+signed(MULTS_3_7(68)(PERCISION) & MULTS_3_7(68)(PERCISION downto 1));
			MULTS_4_4(69)<=signed(MULTS_3_6(69)(PERCISION) & MULTS_3_6(69)(PERCISION downto 1))+signed(MULTS_3_7(69)(PERCISION) & MULTS_3_7(69)(PERCISION downto 1));
			MULTS_4_4(70)<=signed(MULTS_3_6(70)(PERCISION) & MULTS_3_6(70)(PERCISION downto 1))+signed(MULTS_3_7(70)(PERCISION) & MULTS_3_7(70)(PERCISION downto 1));
			MULTS_4_4(71)<=signed(MULTS_3_6(71)(PERCISION) & MULTS_3_6(71)(PERCISION downto 1))+signed(MULTS_3_7(71)(PERCISION) & MULTS_3_7(71)(PERCISION downto 1));
			MULTS_4_4(72)<=signed(MULTS_3_6(72)(PERCISION) & MULTS_3_6(72)(PERCISION downto 1))+signed(MULTS_3_7(72)(PERCISION) & MULTS_3_7(72)(PERCISION downto 1));
			MULTS_4_4(73)<=signed(MULTS_3_6(73)(PERCISION) & MULTS_3_6(73)(PERCISION downto 1))+signed(MULTS_3_7(73)(PERCISION) & MULTS_3_7(73)(PERCISION downto 1));
			MULTS_4_4(74)<=signed(MULTS_3_6(74)(PERCISION) & MULTS_3_6(74)(PERCISION downto 1))+signed(MULTS_3_7(74)(PERCISION) & MULTS_3_7(74)(PERCISION downto 1));
			MULTS_4_4(75)<=signed(MULTS_3_6(75)(PERCISION) & MULTS_3_6(75)(PERCISION downto 1))+signed(MULTS_3_7(75)(PERCISION) & MULTS_3_7(75)(PERCISION downto 1));
			MULTS_4_4(76)<=signed(MULTS_3_6(76)(PERCISION) & MULTS_3_6(76)(PERCISION downto 1))+signed(MULTS_3_7(76)(PERCISION) & MULTS_3_7(76)(PERCISION downto 1));
			MULTS_4_4(77)<=signed(MULTS_3_6(77)(PERCISION) & MULTS_3_6(77)(PERCISION downto 1))+signed(MULTS_3_7(77)(PERCISION) & MULTS_3_7(77)(PERCISION downto 1));
			MULTS_4_4(78)<=signed(MULTS_3_6(78)(PERCISION) & MULTS_3_6(78)(PERCISION downto 1))+signed(MULTS_3_7(78)(PERCISION) & MULTS_3_7(78)(PERCISION downto 1));
			MULTS_4_4(79)<=signed(MULTS_3_6(79)(PERCISION) & MULTS_3_6(79)(PERCISION downto 1))+signed(MULTS_3_7(79)(PERCISION) & MULTS_3_7(79)(PERCISION downto 1));
			MULTS_4_4(80)<=signed(MULTS_3_6(80)(PERCISION) & MULTS_3_6(80)(PERCISION downto 1))+signed(MULTS_3_7(80)(PERCISION) & MULTS_3_7(80)(PERCISION downto 1));
			MULTS_4_4(81)<=signed(MULTS_3_6(81)(PERCISION) & MULTS_3_6(81)(PERCISION downto 1))+signed(MULTS_3_7(81)(PERCISION) & MULTS_3_7(81)(PERCISION downto 1));
			MULTS_4_4(82)<=signed(MULTS_3_6(82)(PERCISION) & MULTS_3_6(82)(PERCISION downto 1))+signed(MULTS_3_7(82)(PERCISION) & MULTS_3_7(82)(PERCISION downto 1));
			MULTS_4_4(83)<=signed(MULTS_3_6(83)(PERCISION) & MULTS_3_6(83)(PERCISION downto 1))+signed(MULTS_3_7(83)(PERCISION) & MULTS_3_7(83)(PERCISION downto 1));

			MULTS_4_5(0)<=signed(MULTS_3_8(0)(PERCISION) & MULTS_3_8(0)(PERCISION downto 1))+signed(MULTS_3_9(0)(PERCISION) & MULTS_3_9(0)(PERCISION downto 1));
			MULTS_4_5(1)<=signed(MULTS_3_8(1)(PERCISION) & MULTS_3_8(1)(PERCISION downto 1))+signed(MULTS_3_9(1)(PERCISION) & MULTS_3_9(1)(PERCISION downto 1));
			MULTS_4_5(2)<=signed(MULTS_3_8(2)(PERCISION) & MULTS_3_8(2)(PERCISION downto 1))+signed(MULTS_3_9(2)(PERCISION) & MULTS_3_9(2)(PERCISION downto 1));
			MULTS_4_5(3)<=signed(MULTS_3_8(3)(PERCISION) & MULTS_3_8(3)(PERCISION downto 1))+signed(MULTS_3_9(3)(PERCISION) & MULTS_3_9(3)(PERCISION downto 1));
			MULTS_4_5(4)<=signed(MULTS_3_8(4)(PERCISION) & MULTS_3_8(4)(PERCISION downto 1))+signed(MULTS_3_9(4)(PERCISION) & MULTS_3_9(4)(PERCISION downto 1));
			MULTS_4_5(5)<=signed(MULTS_3_8(5)(PERCISION) & MULTS_3_8(5)(PERCISION downto 1))+signed(MULTS_3_9(5)(PERCISION) & MULTS_3_9(5)(PERCISION downto 1));
			MULTS_4_5(6)<=signed(MULTS_3_8(6)(PERCISION) & MULTS_3_8(6)(PERCISION downto 1))+signed(MULTS_3_9(6)(PERCISION) & MULTS_3_9(6)(PERCISION downto 1));
			MULTS_4_5(7)<=signed(MULTS_3_8(7)(PERCISION) & MULTS_3_8(7)(PERCISION downto 1))+signed(MULTS_3_9(7)(PERCISION) & MULTS_3_9(7)(PERCISION downto 1));
			MULTS_4_5(8)<=signed(MULTS_3_8(8)(PERCISION) & MULTS_3_8(8)(PERCISION downto 1))+signed(MULTS_3_9(8)(PERCISION) & MULTS_3_9(8)(PERCISION downto 1));
			MULTS_4_5(9)<=signed(MULTS_3_8(9)(PERCISION) & MULTS_3_8(9)(PERCISION downto 1))+signed(MULTS_3_9(9)(PERCISION) & MULTS_3_9(9)(PERCISION downto 1));
			MULTS_4_5(10)<=signed(MULTS_3_8(10)(PERCISION) & MULTS_3_8(10)(PERCISION downto 1))+signed(MULTS_3_9(10)(PERCISION) & MULTS_3_9(10)(PERCISION downto 1));
			MULTS_4_5(11)<=signed(MULTS_3_8(11)(PERCISION) & MULTS_3_8(11)(PERCISION downto 1))+signed(MULTS_3_9(11)(PERCISION) & MULTS_3_9(11)(PERCISION downto 1));
			MULTS_4_5(12)<=signed(MULTS_3_8(12)(PERCISION) & MULTS_3_8(12)(PERCISION downto 1))+signed(MULTS_3_9(12)(PERCISION) & MULTS_3_9(12)(PERCISION downto 1));
			MULTS_4_5(13)<=signed(MULTS_3_8(13)(PERCISION) & MULTS_3_8(13)(PERCISION downto 1))+signed(MULTS_3_9(13)(PERCISION) & MULTS_3_9(13)(PERCISION downto 1));
			MULTS_4_5(14)<=signed(MULTS_3_8(14)(PERCISION) & MULTS_3_8(14)(PERCISION downto 1))+signed(MULTS_3_9(14)(PERCISION) & MULTS_3_9(14)(PERCISION downto 1));
			MULTS_4_5(15)<=signed(MULTS_3_8(15)(PERCISION) & MULTS_3_8(15)(PERCISION downto 1))+signed(MULTS_3_9(15)(PERCISION) & MULTS_3_9(15)(PERCISION downto 1));
			MULTS_4_5(16)<=signed(MULTS_3_8(16)(PERCISION) & MULTS_3_8(16)(PERCISION downto 1))+signed(MULTS_3_9(16)(PERCISION) & MULTS_3_9(16)(PERCISION downto 1));
			MULTS_4_5(17)<=signed(MULTS_3_8(17)(PERCISION) & MULTS_3_8(17)(PERCISION downto 1))+signed(MULTS_3_9(17)(PERCISION) & MULTS_3_9(17)(PERCISION downto 1));
			MULTS_4_5(18)<=signed(MULTS_3_8(18)(PERCISION) & MULTS_3_8(18)(PERCISION downto 1))+signed(MULTS_3_9(18)(PERCISION) & MULTS_3_9(18)(PERCISION downto 1));
			MULTS_4_5(19)<=signed(MULTS_3_8(19)(PERCISION) & MULTS_3_8(19)(PERCISION downto 1))+signed(MULTS_3_9(19)(PERCISION) & MULTS_3_9(19)(PERCISION downto 1));
			MULTS_4_5(20)<=signed(MULTS_3_8(20)(PERCISION) & MULTS_3_8(20)(PERCISION downto 1))+signed(MULTS_3_9(20)(PERCISION) & MULTS_3_9(20)(PERCISION downto 1));
			MULTS_4_5(21)<=signed(MULTS_3_8(21)(PERCISION) & MULTS_3_8(21)(PERCISION downto 1))+signed(MULTS_3_9(21)(PERCISION) & MULTS_3_9(21)(PERCISION downto 1));
			MULTS_4_5(22)<=signed(MULTS_3_8(22)(PERCISION) & MULTS_3_8(22)(PERCISION downto 1))+signed(MULTS_3_9(22)(PERCISION) & MULTS_3_9(22)(PERCISION downto 1));
			MULTS_4_5(23)<=signed(MULTS_3_8(23)(PERCISION) & MULTS_3_8(23)(PERCISION downto 1))+signed(MULTS_3_9(23)(PERCISION) & MULTS_3_9(23)(PERCISION downto 1));
			MULTS_4_5(24)<=signed(MULTS_3_8(24)(PERCISION) & MULTS_3_8(24)(PERCISION downto 1))+signed(MULTS_3_9(24)(PERCISION) & MULTS_3_9(24)(PERCISION downto 1));
			MULTS_4_5(25)<=signed(MULTS_3_8(25)(PERCISION) & MULTS_3_8(25)(PERCISION downto 1))+signed(MULTS_3_9(25)(PERCISION) & MULTS_3_9(25)(PERCISION downto 1));
			MULTS_4_5(26)<=signed(MULTS_3_8(26)(PERCISION) & MULTS_3_8(26)(PERCISION downto 1))+signed(MULTS_3_9(26)(PERCISION) & MULTS_3_9(26)(PERCISION downto 1));
			MULTS_4_5(27)<=signed(MULTS_3_8(27)(PERCISION) & MULTS_3_8(27)(PERCISION downto 1))+signed(MULTS_3_9(27)(PERCISION) & MULTS_3_9(27)(PERCISION downto 1));
			MULTS_4_5(28)<=signed(MULTS_3_8(28)(PERCISION) & MULTS_3_8(28)(PERCISION downto 1))+signed(MULTS_3_9(28)(PERCISION) & MULTS_3_9(28)(PERCISION downto 1));
			MULTS_4_5(29)<=signed(MULTS_3_8(29)(PERCISION) & MULTS_3_8(29)(PERCISION downto 1))+signed(MULTS_3_9(29)(PERCISION) & MULTS_3_9(29)(PERCISION downto 1));
			MULTS_4_5(30)<=signed(MULTS_3_8(30)(PERCISION) & MULTS_3_8(30)(PERCISION downto 1))+signed(MULTS_3_9(30)(PERCISION) & MULTS_3_9(30)(PERCISION downto 1));
			MULTS_4_5(31)<=signed(MULTS_3_8(31)(PERCISION) & MULTS_3_8(31)(PERCISION downto 1))+signed(MULTS_3_9(31)(PERCISION) & MULTS_3_9(31)(PERCISION downto 1));
			MULTS_4_5(32)<=signed(MULTS_3_8(32)(PERCISION) & MULTS_3_8(32)(PERCISION downto 1))+signed(MULTS_3_9(32)(PERCISION) & MULTS_3_9(32)(PERCISION downto 1));
			MULTS_4_5(33)<=signed(MULTS_3_8(33)(PERCISION) & MULTS_3_8(33)(PERCISION downto 1))+signed(MULTS_3_9(33)(PERCISION) & MULTS_3_9(33)(PERCISION downto 1));
			MULTS_4_5(34)<=signed(MULTS_3_8(34)(PERCISION) & MULTS_3_8(34)(PERCISION downto 1))+signed(MULTS_3_9(34)(PERCISION) & MULTS_3_9(34)(PERCISION downto 1));
			MULTS_4_5(35)<=signed(MULTS_3_8(35)(PERCISION) & MULTS_3_8(35)(PERCISION downto 1))+signed(MULTS_3_9(35)(PERCISION) & MULTS_3_9(35)(PERCISION downto 1));
			MULTS_4_5(36)<=signed(MULTS_3_8(36)(PERCISION) & MULTS_3_8(36)(PERCISION downto 1))+signed(MULTS_3_9(36)(PERCISION) & MULTS_3_9(36)(PERCISION downto 1));
			MULTS_4_5(37)<=signed(MULTS_3_8(37)(PERCISION) & MULTS_3_8(37)(PERCISION downto 1))+signed(MULTS_3_9(37)(PERCISION) & MULTS_3_9(37)(PERCISION downto 1));
			MULTS_4_5(38)<=signed(MULTS_3_8(38)(PERCISION) & MULTS_3_8(38)(PERCISION downto 1))+signed(MULTS_3_9(38)(PERCISION) & MULTS_3_9(38)(PERCISION downto 1));
			MULTS_4_5(39)<=signed(MULTS_3_8(39)(PERCISION) & MULTS_3_8(39)(PERCISION downto 1))+signed(MULTS_3_9(39)(PERCISION) & MULTS_3_9(39)(PERCISION downto 1));
			MULTS_4_5(40)<=signed(MULTS_3_8(40)(PERCISION) & MULTS_3_8(40)(PERCISION downto 1))+signed(MULTS_3_9(40)(PERCISION) & MULTS_3_9(40)(PERCISION downto 1));
			MULTS_4_5(41)<=signed(MULTS_3_8(41)(PERCISION) & MULTS_3_8(41)(PERCISION downto 1))+signed(MULTS_3_9(41)(PERCISION) & MULTS_3_9(41)(PERCISION downto 1));
			MULTS_4_5(42)<=signed(MULTS_3_8(42)(PERCISION) & MULTS_3_8(42)(PERCISION downto 1))+signed(MULTS_3_9(42)(PERCISION) & MULTS_3_9(42)(PERCISION downto 1));
			MULTS_4_5(43)<=signed(MULTS_3_8(43)(PERCISION) & MULTS_3_8(43)(PERCISION downto 1))+signed(MULTS_3_9(43)(PERCISION) & MULTS_3_9(43)(PERCISION downto 1));
			MULTS_4_5(44)<=signed(MULTS_3_8(44)(PERCISION) & MULTS_3_8(44)(PERCISION downto 1))+signed(MULTS_3_9(44)(PERCISION) & MULTS_3_9(44)(PERCISION downto 1));
			MULTS_4_5(45)<=signed(MULTS_3_8(45)(PERCISION) & MULTS_3_8(45)(PERCISION downto 1))+signed(MULTS_3_9(45)(PERCISION) & MULTS_3_9(45)(PERCISION downto 1));
			MULTS_4_5(46)<=signed(MULTS_3_8(46)(PERCISION) & MULTS_3_8(46)(PERCISION downto 1))+signed(MULTS_3_9(46)(PERCISION) & MULTS_3_9(46)(PERCISION downto 1));
			MULTS_4_5(47)<=signed(MULTS_3_8(47)(PERCISION) & MULTS_3_8(47)(PERCISION downto 1))+signed(MULTS_3_9(47)(PERCISION) & MULTS_3_9(47)(PERCISION downto 1));
			MULTS_4_5(48)<=signed(MULTS_3_8(48)(PERCISION) & MULTS_3_8(48)(PERCISION downto 1))+signed(MULTS_3_9(48)(PERCISION) & MULTS_3_9(48)(PERCISION downto 1));
			MULTS_4_5(49)<=signed(MULTS_3_8(49)(PERCISION) & MULTS_3_8(49)(PERCISION downto 1))+signed(MULTS_3_9(49)(PERCISION) & MULTS_3_9(49)(PERCISION downto 1));
			MULTS_4_5(50)<=signed(MULTS_3_8(50)(PERCISION) & MULTS_3_8(50)(PERCISION downto 1))+signed(MULTS_3_9(50)(PERCISION) & MULTS_3_9(50)(PERCISION downto 1));
			MULTS_4_5(51)<=signed(MULTS_3_8(51)(PERCISION) & MULTS_3_8(51)(PERCISION downto 1))+signed(MULTS_3_9(51)(PERCISION) & MULTS_3_9(51)(PERCISION downto 1));
			MULTS_4_5(52)<=signed(MULTS_3_8(52)(PERCISION) & MULTS_3_8(52)(PERCISION downto 1))+signed(MULTS_3_9(52)(PERCISION) & MULTS_3_9(52)(PERCISION downto 1));
			MULTS_4_5(53)<=signed(MULTS_3_8(53)(PERCISION) & MULTS_3_8(53)(PERCISION downto 1))+signed(MULTS_3_9(53)(PERCISION) & MULTS_3_9(53)(PERCISION downto 1));
			MULTS_4_5(54)<=signed(MULTS_3_8(54)(PERCISION) & MULTS_3_8(54)(PERCISION downto 1))+signed(MULTS_3_9(54)(PERCISION) & MULTS_3_9(54)(PERCISION downto 1));
			MULTS_4_5(55)<=signed(MULTS_3_8(55)(PERCISION) & MULTS_3_8(55)(PERCISION downto 1))+signed(MULTS_3_9(55)(PERCISION) & MULTS_3_9(55)(PERCISION downto 1));
			MULTS_4_5(56)<=signed(MULTS_3_8(56)(PERCISION) & MULTS_3_8(56)(PERCISION downto 1))+signed(MULTS_3_9(56)(PERCISION) & MULTS_3_9(56)(PERCISION downto 1));
			MULTS_4_5(57)<=signed(MULTS_3_8(57)(PERCISION) & MULTS_3_8(57)(PERCISION downto 1))+signed(MULTS_3_9(57)(PERCISION) & MULTS_3_9(57)(PERCISION downto 1));
			MULTS_4_5(58)<=signed(MULTS_3_8(58)(PERCISION) & MULTS_3_8(58)(PERCISION downto 1))+signed(MULTS_3_9(58)(PERCISION) & MULTS_3_9(58)(PERCISION downto 1));
			MULTS_4_5(59)<=signed(MULTS_3_8(59)(PERCISION) & MULTS_3_8(59)(PERCISION downto 1))+signed(MULTS_3_9(59)(PERCISION) & MULTS_3_9(59)(PERCISION downto 1));
			MULTS_4_5(60)<=signed(MULTS_3_8(60)(PERCISION) & MULTS_3_8(60)(PERCISION downto 1))+signed(MULTS_3_9(60)(PERCISION) & MULTS_3_9(60)(PERCISION downto 1));
			MULTS_4_5(61)<=signed(MULTS_3_8(61)(PERCISION) & MULTS_3_8(61)(PERCISION downto 1))+signed(MULTS_3_9(61)(PERCISION) & MULTS_3_9(61)(PERCISION downto 1));
			MULTS_4_5(62)<=signed(MULTS_3_8(62)(PERCISION) & MULTS_3_8(62)(PERCISION downto 1))+signed(MULTS_3_9(62)(PERCISION) & MULTS_3_9(62)(PERCISION downto 1));
			MULTS_4_5(63)<=signed(MULTS_3_8(63)(PERCISION) & MULTS_3_8(63)(PERCISION downto 1))+signed(MULTS_3_9(63)(PERCISION) & MULTS_3_9(63)(PERCISION downto 1));
			MULTS_4_5(64)<=signed(MULTS_3_8(64)(PERCISION) & MULTS_3_8(64)(PERCISION downto 1))+signed(MULTS_3_9(64)(PERCISION) & MULTS_3_9(64)(PERCISION downto 1));
			MULTS_4_5(65)<=signed(MULTS_3_8(65)(PERCISION) & MULTS_3_8(65)(PERCISION downto 1))+signed(MULTS_3_9(65)(PERCISION) & MULTS_3_9(65)(PERCISION downto 1));
			MULTS_4_5(66)<=signed(MULTS_3_8(66)(PERCISION) & MULTS_3_8(66)(PERCISION downto 1))+signed(MULTS_3_9(66)(PERCISION) & MULTS_3_9(66)(PERCISION downto 1));
			MULTS_4_5(67)<=signed(MULTS_3_8(67)(PERCISION) & MULTS_3_8(67)(PERCISION downto 1))+signed(MULTS_3_9(67)(PERCISION) & MULTS_3_9(67)(PERCISION downto 1));
			MULTS_4_5(68)<=signed(MULTS_3_8(68)(PERCISION) & MULTS_3_8(68)(PERCISION downto 1))+signed(MULTS_3_9(68)(PERCISION) & MULTS_3_9(68)(PERCISION downto 1));
			MULTS_4_5(69)<=signed(MULTS_3_8(69)(PERCISION) & MULTS_3_8(69)(PERCISION downto 1))+signed(MULTS_3_9(69)(PERCISION) & MULTS_3_9(69)(PERCISION downto 1));
			MULTS_4_5(70)<=signed(MULTS_3_8(70)(PERCISION) & MULTS_3_8(70)(PERCISION downto 1))+signed(MULTS_3_9(70)(PERCISION) & MULTS_3_9(70)(PERCISION downto 1));
			MULTS_4_5(71)<=signed(MULTS_3_8(71)(PERCISION) & MULTS_3_8(71)(PERCISION downto 1))+signed(MULTS_3_9(71)(PERCISION) & MULTS_3_9(71)(PERCISION downto 1));
			MULTS_4_5(72)<=signed(MULTS_3_8(72)(PERCISION) & MULTS_3_8(72)(PERCISION downto 1))+signed(MULTS_3_9(72)(PERCISION) & MULTS_3_9(72)(PERCISION downto 1));
			MULTS_4_5(73)<=signed(MULTS_3_8(73)(PERCISION) & MULTS_3_8(73)(PERCISION downto 1))+signed(MULTS_3_9(73)(PERCISION) & MULTS_3_9(73)(PERCISION downto 1));
			MULTS_4_5(74)<=signed(MULTS_3_8(74)(PERCISION) & MULTS_3_8(74)(PERCISION downto 1))+signed(MULTS_3_9(74)(PERCISION) & MULTS_3_9(74)(PERCISION downto 1));
			MULTS_4_5(75)<=signed(MULTS_3_8(75)(PERCISION) & MULTS_3_8(75)(PERCISION downto 1))+signed(MULTS_3_9(75)(PERCISION) & MULTS_3_9(75)(PERCISION downto 1));
			MULTS_4_5(76)<=signed(MULTS_3_8(76)(PERCISION) & MULTS_3_8(76)(PERCISION downto 1))+signed(MULTS_3_9(76)(PERCISION) & MULTS_3_9(76)(PERCISION downto 1));
			MULTS_4_5(77)<=signed(MULTS_3_8(77)(PERCISION) & MULTS_3_8(77)(PERCISION downto 1))+signed(MULTS_3_9(77)(PERCISION) & MULTS_3_9(77)(PERCISION downto 1));
			MULTS_4_5(78)<=signed(MULTS_3_8(78)(PERCISION) & MULTS_3_8(78)(PERCISION downto 1))+signed(MULTS_3_9(78)(PERCISION) & MULTS_3_9(78)(PERCISION downto 1));
			MULTS_4_5(79)<=signed(MULTS_3_8(79)(PERCISION) & MULTS_3_8(79)(PERCISION downto 1))+signed(MULTS_3_9(79)(PERCISION) & MULTS_3_9(79)(PERCISION downto 1));
			MULTS_4_5(80)<=signed(MULTS_3_8(80)(PERCISION) & MULTS_3_8(80)(PERCISION downto 1))+signed(MULTS_3_9(80)(PERCISION) & MULTS_3_9(80)(PERCISION downto 1));
			MULTS_4_5(81)<=signed(MULTS_3_8(81)(PERCISION) & MULTS_3_8(81)(PERCISION downto 1))+signed(MULTS_3_9(81)(PERCISION) & MULTS_3_9(81)(PERCISION downto 1));
			MULTS_4_5(82)<=signed(MULTS_3_8(82)(PERCISION) & MULTS_3_8(82)(PERCISION downto 1))+signed(MULTS_3_9(82)(PERCISION) & MULTS_3_9(82)(PERCISION downto 1));
			MULTS_4_5(83)<=signed(MULTS_3_8(83)(PERCISION) & MULTS_3_8(83)(PERCISION downto 1))+signed(MULTS_3_9(83)(PERCISION) & MULTS_3_9(83)(PERCISION downto 1));



                         EN_SUM_MULT_5<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_5 = '1' then
			------------------------------------STAGE-5--------------------------------------
			MULTS_5_1(0)<=signed(MULTS_4_1(0)(PERCISION) & MULTS_4_1(0)(PERCISION downto 1))+signed(MULTS_4_2(0)(PERCISION) & MULTS_4_2(0)(PERCISION downto 1));
			MULTS_5_1(1)<=signed(MULTS_4_1(1)(PERCISION) & MULTS_4_1(1)(PERCISION downto 1))+signed(MULTS_4_2(1)(PERCISION) & MULTS_4_2(1)(PERCISION downto 1));
			MULTS_5_1(2)<=signed(MULTS_4_1(2)(PERCISION) & MULTS_4_1(2)(PERCISION downto 1))+signed(MULTS_4_2(2)(PERCISION) & MULTS_4_2(2)(PERCISION downto 1));
			MULTS_5_1(3)<=signed(MULTS_4_1(3)(PERCISION) & MULTS_4_1(3)(PERCISION downto 1))+signed(MULTS_4_2(3)(PERCISION) & MULTS_4_2(3)(PERCISION downto 1));
			MULTS_5_1(4)<=signed(MULTS_4_1(4)(PERCISION) & MULTS_4_1(4)(PERCISION downto 1))+signed(MULTS_4_2(4)(PERCISION) & MULTS_4_2(4)(PERCISION downto 1));
			MULTS_5_1(5)<=signed(MULTS_4_1(5)(PERCISION) & MULTS_4_1(5)(PERCISION downto 1))+signed(MULTS_4_2(5)(PERCISION) & MULTS_4_2(5)(PERCISION downto 1));
			MULTS_5_1(6)<=signed(MULTS_4_1(6)(PERCISION) & MULTS_4_1(6)(PERCISION downto 1))+signed(MULTS_4_2(6)(PERCISION) & MULTS_4_2(6)(PERCISION downto 1));
			MULTS_5_1(7)<=signed(MULTS_4_1(7)(PERCISION) & MULTS_4_1(7)(PERCISION downto 1))+signed(MULTS_4_2(7)(PERCISION) & MULTS_4_2(7)(PERCISION downto 1));
			MULTS_5_1(8)<=signed(MULTS_4_1(8)(PERCISION) & MULTS_4_1(8)(PERCISION downto 1))+signed(MULTS_4_2(8)(PERCISION) & MULTS_4_2(8)(PERCISION downto 1));
			MULTS_5_1(9)<=signed(MULTS_4_1(9)(PERCISION) & MULTS_4_1(9)(PERCISION downto 1))+signed(MULTS_4_2(9)(PERCISION) & MULTS_4_2(9)(PERCISION downto 1));
			MULTS_5_1(10)<=signed(MULTS_4_1(10)(PERCISION) & MULTS_4_1(10)(PERCISION downto 1))+signed(MULTS_4_2(10)(PERCISION) & MULTS_4_2(10)(PERCISION downto 1));
			MULTS_5_1(11)<=signed(MULTS_4_1(11)(PERCISION) & MULTS_4_1(11)(PERCISION downto 1))+signed(MULTS_4_2(11)(PERCISION) & MULTS_4_2(11)(PERCISION downto 1));
			MULTS_5_1(12)<=signed(MULTS_4_1(12)(PERCISION) & MULTS_4_1(12)(PERCISION downto 1))+signed(MULTS_4_2(12)(PERCISION) & MULTS_4_2(12)(PERCISION downto 1));
			MULTS_5_1(13)<=signed(MULTS_4_1(13)(PERCISION) & MULTS_4_1(13)(PERCISION downto 1))+signed(MULTS_4_2(13)(PERCISION) & MULTS_4_2(13)(PERCISION downto 1));
			MULTS_5_1(14)<=signed(MULTS_4_1(14)(PERCISION) & MULTS_4_1(14)(PERCISION downto 1))+signed(MULTS_4_2(14)(PERCISION) & MULTS_4_2(14)(PERCISION downto 1));
			MULTS_5_1(15)<=signed(MULTS_4_1(15)(PERCISION) & MULTS_4_1(15)(PERCISION downto 1))+signed(MULTS_4_2(15)(PERCISION) & MULTS_4_2(15)(PERCISION downto 1));
			MULTS_5_1(16)<=signed(MULTS_4_1(16)(PERCISION) & MULTS_4_1(16)(PERCISION downto 1))+signed(MULTS_4_2(16)(PERCISION) & MULTS_4_2(16)(PERCISION downto 1));
			MULTS_5_1(17)<=signed(MULTS_4_1(17)(PERCISION) & MULTS_4_1(17)(PERCISION downto 1))+signed(MULTS_4_2(17)(PERCISION) & MULTS_4_2(17)(PERCISION downto 1));
			MULTS_5_1(18)<=signed(MULTS_4_1(18)(PERCISION) & MULTS_4_1(18)(PERCISION downto 1))+signed(MULTS_4_2(18)(PERCISION) & MULTS_4_2(18)(PERCISION downto 1));
			MULTS_5_1(19)<=signed(MULTS_4_1(19)(PERCISION) & MULTS_4_1(19)(PERCISION downto 1))+signed(MULTS_4_2(19)(PERCISION) & MULTS_4_2(19)(PERCISION downto 1));
			MULTS_5_1(20)<=signed(MULTS_4_1(20)(PERCISION) & MULTS_4_1(20)(PERCISION downto 1))+signed(MULTS_4_2(20)(PERCISION) & MULTS_4_2(20)(PERCISION downto 1));
			MULTS_5_1(21)<=signed(MULTS_4_1(21)(PERCISION) & MULTS_4_1(21)(PERCISION downto 1))+signed(MULTS_4_2(21)(PERCISION) & MULTS_4_2(21)(PERCISION downto 1));
			MULTS_5_1(22)<=signed(MULTS_4_1(22)(PERCISION) & MULTS_4_1(22)(PERCISION downto 1))+signed(MULTS_4_2(22)(PERCISION) & MULTS_4_2(22)(PERCISION downto 1));
			MULTS_5_1(23)<=signed(MULTS_4_1(23)(PERCISION) & MULTS_4_1(23)(PERCISION downto 1))+signed(MULTS_4_2(23)(PERCISION) & MULTS_4_2(23)(PERCISION downto 1));
			MULTS_5_1(24)<=signed(MULTS_4_1(24)(PERCISION) & MULTS_4_1(24)(PERCISION downto 1))+signed(MULTS_4_2(24)(PERCISION) & MULTS_4_2(24)(PERCISION downto 1));
			MULTS_5_1(25)<=signed(MULTS_4_1(25)(PERCISION) & MULTS_4_1(25)(PERCISION downto 1))+signed(MULTS_4_2(25)(PERCISION) & MULTS_4_2(25)(PERCISION downto 1));
			MULTS_5_1(26)<=signed(MULTS_4_1(26)(PERCISION) & MULTS_4_1(26)(PERCISION downto 1))+signed(MULTS_4_2(26)(PERCISION) & MULTS_4_2(26)(PERCISION downto 1));
			MULTS_5_1(27)<=signed(MULTS_4_1(27)(PERCISION) & MULTS_4_1(27)(PERCISION downto 1))+signed(MULTS_4_2(27)(PERCISION) & MULTS_4_2(27)(PERCISION downto 1));
			MULTS_5_1(28)<=signed(MULTS_4_1(28)(PERCISION) & MULTS_4_1(28)(PERCISION downto 1))+signed(MULTS_4_2(28)(PERCISION) & MULTS_4_2(28)(PERCISION downto 1));
			MULTS_5_1(29)<=signed(MULTS_4_1(29)(PERCISION) & MULTS_4_1(29)(PERCISION downto 1))+signed(MULTS_4_2(29)(PERCISION) & MULTS_4_2(29)(PERCISION downto 1));
			MULTS_5_1(30)<=signed(MULTS_4_1(30)(PERCISION) & MULTS_4_1(30)(PERCISION downto 1))+signed(MULTS_4_2(30)(PERCISION) & MULTS_4_2(30)(PERCISION downto 1));
			MULTS_5_1(31)<=signed(MULTS_4_1(31)(PERCISION) & MULTS_4_1(31)(PERCISION downto 1))+signed(MULTS_4_2(31)(PERCISION) & MULTS_4_2(31)(PERCISION downto 1));
			MULTS_5_1(32)<=signed(MULTS_4_1(32)(PERCISION) & MULTS_4_1(32)(PERCISION downto 1))+signed(MULTS_4_2(32)(PERCISION) & MULTS_4_2(32)(PERCISION downto 1));
			MULTS_5_1(33)<=signed(MULTS_4_1(33)(PERCISION) & MULTS_4_1(33)(PERCISION downto 1))+signed(MULTS_4_2(33)(PERCISION) & MULTS_4_2(33)(PERCISION downto 1));
			MULTS_5_1(34)<=signed(MULTS_4_1(34)(PERCISION) & MULTS_4_1(34)(PERCISION downto 1))+signed(MULTS_4_2(34)(PERCISION) & MULTS_4_2(34)(PERCISION downto 1));
			MULTS_5_1(35)<=signed(MULTS_4_1(35)(PERCISION) & MULTS_4_1(35)(PERCISION downto 1))+signed(MULTS_4_2(35)(PERCISION) & MULTS_4_2(35)(PERCISION downto 1));
			MULTS_5_1(36)<=signed(MULTS_4_1(36)(PERCISION) & MULTS_4_1(36)(PERCISION downto 1))+signed(MULTS_4_2(36)(PERCISION) & MULTS_4_2(36)(PERCISION downto 1));
			MULTS_5_1(37)<=signed(MULTS_4_1(37)(PERCISION) & MULTS_4_1(37)(PERCISION downto 1))+signed(MULTS_4_2(37)(PERCISION) & MULTS_4_2(37)(PERCISION downto 1));
			MULTS_5_1(38)<=signed(MULTS_4_1(38)(PERCISION) & MULTS_4_1(38)(PERCISION downto 1))+signed(MULTS_4_2(38)(PERCISION) & MULTS_4_2(38)(PERCISION downto 1));
			MULTS_5_1(39)<=signed(MULTS_4_1(39)(PERCISION) & MULTS_4_1(39)(PERCISION downto 1))+signed(MULTS_4_2(39)(PERCISION) & MULTS_4_2(39)(PERCISION downto 1));
			MULTS_5_1(40)<=signed(MULTS_4_1(40)(PERCISION) & MULTS_4_1(40)(PERCISION downto 1))+signed(MULTS_4_2(40)(PERCISION) & MULTS_4_2(40)(PERCISION downto 1));
			MULTS_5_1(41)<=signed(MULTS_4_1(41)(PERCISION) & MULTS_4_1(41)(PERCISION downto 1))+signed(MULTS_4_2(41)(PERCISION) & MULTS_4_2(41)(PERCISION downto 1));
			MULTS_5_1(42)<=signed(MULTS_4_1(42)(PERCISION) & MULTS_4_1(42)(PERCISION downto 1))+signed(MULTS_4_2(42)(PERCISION) & MULTS_4_2(42)(PERCISION downto 1));
			MULTS_5_1(43)<=signed(MULTS_4_1(43)(PERCISION) & MULTS_4_1(43)(PERCISION downto 1))+signed(MULTS_4_2(43)(PERCISION) & MULTS_4_2(43)(PERCISION downto 1));
			MULTS_5_1(44)<=signed(MULTS_4_1(44)(PERCISION) & MULTS_4_1(44)(PERCISION downto 1))+signed(MULTS_4_2(44)(PERCISION) & MULTS_4_2(44)(PERCISION downto 1));
			MULTS_5_1(45)<=signed(MULTS_4_1(45)(PERCISION) & MULTS_4_1(45)(PERCISION downto 1))+signed(MULTS_4_2(45)(PERCISION) & MULTS_4_2(45)(PERCISION downto 1));
			MULTS_5_1(46)<=signed(MULTS_4_1(46)(PERCISION) & MULTS_4_1(46)(PERCISION downto 1))+signed(MULTS_4_2(46)(PERCISION) & MULTS_4_2(46)(PERCISION downto 1));
			MULTS_5_1(47)<=signed(MULTS_4_1(47)(PERCISION) & MULTS_4_1(47)(PERCISION downto 1))+signed(MULTS_4_2(47)(PERCISION) & MULTS_4_2(47)(PERCISION downto 1));
			MULTS_5_1(48)<=signed(MULTS_4_1(48)(PERCISION) & MULTS_4_1(48)(PERCISION downto 1))+signed(MULTS_4_2(48)(PERCISION) & MULTS_4_2(48)(PERCISION downto 1));
			MULTS_5_1(49)<=signed(MULTS_4_1(49)(PERCISION) & MULTS_4_1(49)(PERCISION downto 1))+signed(MULTS_4_2(49)(PERCISION) & MULTS_4_2(49)(PERCISION downto 1));
			MULTS_5_1(50)<=signed(MULTS_4_1(50)(PERCISION) & MULTS_4_1(50)(PERCISION downto 1))+signed(MULTS_4_2(50)(PERCISION) & MULTS_4_2(50)(PERCISION downto 1));
			MULTS_5_1(51)<=signed(MULTS_4_1(51)(PERCISION) & MULTS_4_1(51)(PERCISION downto 1))+signed(MULTS_4_2(51)(PERCISION) & MULTS_4_2(51)(PERCISION downto 1));
			MULTS_5_1(52)<=signed(MULTS_4_1(52)(PERCISION) & MULTS_4_1(52)(PERCISION downto 1))+signed(MULTS_4_2(52)(PERCISION) & MULTS_4_2(52)(PERCISION downto 1));
			MULTS_5_1(53)<=signed(MULTS_4_1(53)(PERCISION) & MULTS_4_1(53)(PERCISION downto 1))+signed(MULTS_4_2(53)(PERCISION) & MULTS_4_2(53)(PERCISION downto 1));
			MULTS_5_1(54)<=signed(MULTS_4_1(54)(PERCISION) & MULTS_4_1(54)(PERCISION downto 1))+signed(MULTS_4_2(54)(PERCISION) & MULTS_4_2(54)(PERCISION downto 1));
			MULTS_5_1(55)<=signed(MULTS_4_1(55)(PERCISION) & MULTS_4_1(55)(PERCISION downto 1))+signed(MULTS_4_2(55)(PERCISION) & MULTS_4_2(55)(PERCISION downto 1));
			MULTS_5_1(56)<=signed(MULTS_4_1(56)(PERCISION) & MULTS_4_1(56)(PERCISION downto 1))+signed(MULTS_4_2(56)(PERCISION) & MULTS_4_2(56)(PERCISION downto 1));
			MULTS_5_1(57)<=signed(MULTS_4_1(57)(PERCISION) & MULTS_4_1(57)(PERCISION downto 1))+signed(MULTS_4_2(57)(PERCISION) & MULTS_4_2(57)(PERCISION downto 1));
			MULTS_5_1(58)<=signed(MULTS_4_1(58)(PERCISION) & MULTS_4_1(58)(PERCISION downto 1))+signed(MULTS_4_2(58)(PERCISION) & MULTS_4_2(58)(PERCISION downto 1));
			MULTS_5_1(59)<=signed(MULTS_4_1(59)(PERCISION) & MULTS_4_1(59)(PERCISION downto 1))+signed(MULTS_4_2(59)(PERCISION) & MULTS_4_2(59)(PERCISION downto 1));
			MULTS_5_1(60)<=signed(MULTS_4_1(60)(PERCISION) & MULTS_4_1(60)(PERCISION downto 1))+signed(MULTS_4_2(60)(PERCISION) & MULTS_4_2(60)(PERCISION downto 1));
			MULTS_5_1(61)<=signed(MULTS_4_1(61)(PERCISION) & MULTS_4_1(61)(PERCISION downto 1))+signed(MULTS_4_2(61)(PERCISION) & MULTS_4_2(61)(PERCISION downto 1));
			MULTS_5_1(62)<=signed(MULTS_4_1(62)(PERCISION) & MULTS_4_1(62)(PERCISION downto 1))+signed(MULTS_4_2(62)(PERCISION) & MULTS_4_2(62)(PERCISION downto 1));
			MULTS_5_1(63)<=signed(MULTS_4_1(63)(PERCISION) & MULTS_4_1(63)(PERCISION downto 1))+signed(MULTS_4_2(63)(PERCISION) & MULTS_4_2(63)(PERCISION downto 1));
			MULTS_5_1(64)<=signed(MULTS_4_1(64)(PERCISION) & MULTS_4_1(64)(PERCISION downto 1))+signed(MULTS_4_2(64)(PERCISION) & MULTS_4_2(64)(PERCISION downto 1));
			MULTS_5_1(65)<=signed(MULTS_4_1(65)(PERCISION) & MULTS_4_1(65)(PERCISION downto 1))+signed(MULTS_4_2(65)(PERCISION) & MULTS_4_2(65)(PERCISION downto 1));
			MULTS_5_1(66)<=signed(MULTS_4_1(66)(PERCISION) & MULTS_4_1(66)(PERCISION downto 1))+signed(MULTS_4_2(66)(PERCISION) & MULTS_4_2(66)(PERCISION downto 1));
			MULTS_5_1(67)<=signed(MULTS_4_1(67)(PERCISION) & MULTS_4_1(67)(PERCISION downto 1))+signed(MULTS_4_2(67)(PERCISION) & MULTS_4_2(67)(PERCISION downto 1));
			MULTS_5_1(68)<=signed(MULTS_4_1(68)(PERCISION) & MULTS_4_1(68)(PERCISION downto 1))+signed(MULTS_4_2(68)(PERCISION) & MULTS_4_2(68)(PERCISION downto 1));
			MULTS_5_1(69)<=signed(MULTS_4_1(69)(PERCISION) & MULTS_4_1(69)(PERCISION downto 1))+signed(MULTS_4_2(69)(PERCISION) & MULTS_4_2(69)(PERCISION downto 1));
			MULTS_5_1(70)<=signed(MULTS_4_1(70)(PERCISION) & MULTS_4_1(70)(PERCISION downto 1))+signed(MULTS_4_2(70)(PERCISION) & MULTS_4_2(70)(PERCISION downto 1));
			MULTS_5_1(71)<=signed(MULTS_4_1(71)(PERCISION) & MULTS_4_1(71)(PERCISION downto 1))+signed(MULTS_4_2(71)(PERCISION) & MULTS_4_2(71)(PERCISION downto 1));
			MULTS_5_1(72)<=signed(MULTS_4_1(72)(PERCISION) & MULTS_4_1(72)(PERCISION downto 1))+signed(MULTS_4_2(72)(PERCISION) & MULTS_4_2(72)(PERCISION downto 1));
			MULTS_5_1(73)<=signed(MULTS_4_1(73)(PERCISION) & MULTS_4_1(73)(PERCISION downto 1))+signed(MULTS_4_2(73)(PERCISION) & MULTS_4_2(73)(PERCISION downto 1));
			MULTS_5_1(74)<=signed(MULTS_4_1(74)(PERCISION) & MULTS_4_1(74)(PERCISION downto 1))+signed(MULTS_4_2(74)(PERCISION) & MULTS_4_2(74)(PERCISION downto 1));
			MULTS_5_1(75)<=signed(MULTS_4_1(75)(PERCISION) & MULTS_4_1(75)(PERCISION downto 1))+signed(MULTS_4_2(75)(PERCISION) & MULTS_4_2(75)(PERCISION downto 1));
			MULTS_5_1(76)<=signed(MULTS_4_1(76)(PERCISION) & MULTS_4_1(76)(PERCISION downto 1))+signed(MULTS_4_2(76)(PERCISION) & MULTS_4_2(76)(PERCISION downto 1));
			MULTS_5_1(77)<=signed(MULTS_4_1(77)(PERCISION) & MULTS_4_1(77)(PERCISION downto 1))+signed(MULTS_4_2(77)(PERCISION) & MULTS_4_2(77)(PERCISION downto 1));
			MULTS_5_1(78)<=signed(MULTS_4_1(78)(PERCISION) & MULTS_4_1(78)(PERCISION downto 1))+signed(MULTS_4_2(78)(PERCISION) & MULTS_4_2(78)(PERCISION downto 1));
			MULTS_5_1(79)<=signed(MULTS_4_1(79)(PERCISION) & MULTS_4_1(79)(PERCISION downto 1))+signed(MULTS_4_2(79)(PERCISION) & MULTS_4_2(79)(PERCISION downto 1));
			MULTS_5_1(80)<=signed(MULTS_4_1(80)(PERCISION) & MULTS_4_1(80)(PERCISION downto 1))+signed(MULTS_4_2(80)(PERCISION) & MULTS_4_2(80)(PERCISION downto 1));
			MULTS_5_1(81)<=signed(MULTS_4_1(81)(PERCISION) & MULTS_4_1(81)(PERCISION downto 1))+signed(MULTS_4_2(81)(PERCISION) & MULTS_4_2(81)(PERCISION downto 1));
			MULTS_5_1(82)<=signed(MULTS_4_1(82)(PERCISION) & MULTS_4_1(82)(PERCISION downto 1))+signed(MULTS_4_2(82)(PERCISION) & MULTS_4_2(82)(PERCISION downto 1));
			MULTS_5_1(83)<=signed(MULTS_4_1(83)(PERCISION) & MULTS_4_1(83)(PERCISION downto 1))+signed(MULTS_4_2(83)(PERCISION) & MULTS_4_2(83)(PERCISION downto 1));

			MULTS_5_2(0)<=signed(MULTS_4_3(0)(PERCISION) & MULTS_4_3(0)(PERCISION downto 1))+signed(MULTS_4_4(0)(PERCISION) & MULTS_4_4(0)(PERCISION downto 1));
			MULTS_5_2(1)<=signed(MULTS_4_3(1)(PERCISION) & MULTS_4_3(1)(PERCISION downto 1))+signed(MULTS_4_4(1)(PERCISION) & MULTS_4_4(1)(PERCISION downto 1));
			MULTS_5_2(2)<=signed(MULTS_4_3(2)(PERCISION) & MULTS_4_3(2)(PERCISION downto 1))+signed(MULTS_4_4(2)(PERCISION) & MULTS_4_4(2)(PERCISION downto 1));
			MULTS_5_2(3)<=signed(MULTS_4_3(3)(PERCISION) & MULTS_4_3(3)(PERCISION downto 1))+signed(MULTS_4_4(3)(PERCISION) & MULTS_4_4(3)(PERCISION downto 1));
			MULTS_5_2(4)<=signed(MULTS_4_3(4)(PERCISION) & MULTS_4_3(4)(PERCISION downto 1))+signed(MULTS_4_4(4)(PERCISION) & MULTS_4_4(4)(PERCISION downto 1));
			MULTS_5_2(5)<=signed(MULTS_4_3(5)(PERCISION) & MULTS_4_3(5)(PERCISION downto 1))+signed(MULTS_4_4(5)(PERCISION) & MULTS_4_4(5)(PERCISION downto 1));
			MULTS_5_2(6)<=signed(MULTS_4_3(6)(PERCISION) & MULTS_4_3(6)(PERCISION downto 1))+signed(MULTS_4_4(6)(PERCISION) & MULTS_4_4(6)(PERCISION downto 1));
			MULTS_5_2(7)<=signed(MULTS_4_3(7)(PERCISION) & MULTS_4_3(7)(PERCISION downto 1))+signed(MULTS_4_4(7)(PERCISION) & MULTS_4_4(7)(PERCISION downto 1));
			MULTS_5_2(8)<=signed(MULTS_4_3(8)(PERCISION) & MULTS_4_3(8)(PERCISION downto 1))+signed(MULTS_4_4(8)(PERCISION) & MULTS_4_4(8)(PERCISION downto 1));
			MULTS_5_2(9)<=signed(MULTS_4_3(9)(PERCISION) & MULTS_4_3(9)(PERCISION downto 1))+signed(MULTS_4_4(9)(PERCISION) & MULTS_4_4(9)(PERCISION downto 1));
			MULTS_5_2(10)<=signed(MULTS_4_3(10)(PERCISION) & MULTS_4_3(10)(PERCISION downto 1))+signed(MULTS_4_4(10)(PERCISION) & MULTS_4_4(10)(PERCISION downto 1));
			MULTS_5_2(11)<=signed(MULTS_4_3(11)(PERCISION) & MULTS_4_3(11)(PERCISION downto 1))+signed(MULTS_4_4(11)(PERCISION) & MULTS_4_4(11)(PERCISION downto 1));
			MULTS_5_2(12)<=signed(MULTS_4_3(12)(PERCISION) & MULTS_4_3(12)(PERCISION downto 1))+signed(MULTS_4_4(12)(PERCISION) & MULTS_4_4(12)(PERCISION downto 1));
			MULTS_5_2(13)<=signed(MULTS_4_3(13)(PERCISION) & MULTS_4_3(13)(PERCISION downto 1))+signed(MULTS_4_4(13)(PERCISION) & MULTS_4_4(13)(PERCISION downto 1));
			MULTS_5_2(14)<=signed(MULTS_4_3(14)(PERCISION) & MULTS_4_3(14)(PERCISION downto 1))+signed(MULTS_4_4(14)(PERCISION) & MULTS_4_4(14)(PERCISION downto 1));
			MULTS_5_2(15)<=signed(MULTS_4_3(15)(PERCISION) & MULTS_4_3(15)(PERCISION downto 1))+signed(MULTS_4_4(15)(PERCISION) & MULTS_4_4(15)(PERCISION downto 1));
			MULTS_5_2(16)<=signed(MULTS_4_3(16)(PERCISION) & MULTS_4_3(16)(PERCISION downto 1))+signed(MULTS_4_4(16)(PERCISION) & MULTS_4_4(16)(PERCISION downto 1));
			MULTS_5_2(17)<=signed(MULTS_4_3(17)(PERCISION) & MULTS_4_3(17)(PERCISION downto 1))+signed(MULTS_4_4(17)(PERCISION) & MULTS_4_4(17)(PERCISION downto 1));
			MULTS_5_2(18)<=signed(MULTS_4_3(18)(PERCISION) & MULTS_4_3(18)(PERCISION downto 1))+signed(MULTS_4_4(18)(PERCISION) & MULTS_4_4(18)(PERCISION downto 1));
			MULTS_5_2(19)<=signed(MULTS_4_3(19)(PERCISION) & MULTS_4_3(19)(PERCISION downto 1))+signed(MULTS_4_4(19)(PERCISION) & MULTS_4_4(19)(PERCISION downto 1));
			MULTS_5_2(20)<=signed(MULTS_4_3(20)(PERCISION) & MULTS_4_3(20)(PERCISION downto 1))+signed(MULTS_4_4(20)(PERCISION) & MULTS_4_4(20)(PERCISION downto 1));
			MULTS_5_2(21)<=signed(MULTS_4_3(21)(PERCISION) & MULTS_4_3(21)(PERCISION downto 1))+signed(MULTS_4_4(21)(PERCISION) & MULTS_4_4(21)(PERCISION downto 1));
			MULTS_5_2(22)<=signed(MULTS_4_3(22)(PERCISION) & MULTS_4_3(22)(PERCISION downto 1))+signed(MULTS_4_4(22)(PERCISION) & MULTS_4_4(22)(PERCISION downto 1));
			MULTS_5_2(23)<=signed(MULTS_4_3(23)(PERCISION) & MULTS_4_3(23)(PERCISION downto 1))+signed(MULTS_4_4(23)(PERCISION) & MULTS_4_4(23)(PERCISION downto 1));
			MULTS_5_2(24)<=signed(MULTS_4_3(24)(PERCISION) & MULTS_4_3(24)(PERCISION downto 1))+signed(MULTS_4_4(24)(PERCISION) & MULTS_4_4(24)(PERCISION downto 1));
			MULTS_5_2(25)<=signed(MULTS_4_3(25)(PERCISION) & MULTS_4_3(25)(PERCISION downto 1))+signed(MULTS_4_4(25)(PERCISION) & MULTS_4_4(25)(PERCISION downto 1));
			MULTS_5_2(26)<=signed(MULTS_4_3(26)(PERCISION) & MULTS_4_3(26)(PERCISION downto 1))+signed(MULTS_4_4(26)(PERCISION) & MULTS_4_4(26)(PERCISION downto 1));
			MULTS_5_2(27)<=signed(MULTS_4_3(27)(PERCISION) & MULTS_4_3(27)(PERCISION downto 1))+signed(MULTS_4_4(27)(PERCISION) & MULTS_4_4(27)(PERCISION downto 1));
			MULTS_5_2(28)<=signed(MULTS_4_3(28)(PERCISION) & MULTS_4_3(28)(PERCISION downto 1))+signed(MULTS_4_4(28)(PERCISION) & MULTS_4_4(28)(PERCISION downto 1));
			MULTS_5_2(29)<=signed(MULTS_4_3(29)(PERCISION) & MULTS_4_3(29)(PERCISION downto 1))+signed(MULTS_4_4(29)(PERCISION) & MULTS_4_4(29)(PERCISION downto 1));
			MULTS_5_2(30)<=signed(MULTS_4_3(30)(PERCISION) & MULTS_4_3(30)(PERCISION downto 1))+signed(MULTS_4_4(30)(PERCISION) & MULTS_4_4(30)(PERCISION downto 1));
			MULTS_5_2(31)<=signed(MULTS_4_3(31)(PERCISION) & MULTS_4_3(31)(PERCISION downto 1))+signed(MULTS_4_4(31)(PERCISION) & MULTS_4_4(31)(PERCISION downto 1));
			MULTS_5_2(32)<=signed(MULTS_4_3(32)(PERCISION) & MULTS_4_3(32)(PERCISION downto 1))+signed(MULTS_4_4(32)(PERCISION) & MULTS_4_4(32)(PERCISION downto 1));
			MULTS_5_2(33)<=signed(MULTS_4_3(33)(PERCISION) & MULTS_4_3(33)(PERCISION downto 1))+signed(MULTS_4_4(33)(PERCISION) & MULTS_4_4(33)(PERCISION downto 1));
			MULTS_5_2(34)<=signed(MULTS_4_3(34)(PERCISION) & MULTS_4_3(34)(PERCISION downto 1))+signed(MULTS_4_4(34)(PERCISION) & MULTS_4_4(34)(PERCISION downto 1));
			MULTS_5_2(35)<=signed(MULTS_4_3(35)(PERCISION) & MULTS_4_3(35)(PERCISION downto 1))+signed(MULTS_4_4(35)(PERCISION) & MULTS_4_4(35)(PERCISION downto 1));
			MULTS_5_2(36)<=signed(MULTS_4_3(36)(PERCISION) & MULTS_4_3(36)(PERCISION downto 1))+signed(MULTS_4_4(36)(PERCISION) & MULTS_4_4(36)(PERCISION downto 1));
			MULTS_5_2(37)<=signed(MULTS_4_3(37)(PERCISION) & MULTS_4_3(37)(PERCISION downto 1))+signed(MULTS_4_4(37)(PERCISION) & MULTS_4_4(37)(PERCISION downto 1));
			MULTS_5_2(38)<=signed(MULTS_4_3(38)(PERCISION) & MULTS_4_3(38)(PERCISION downto 1))+signed(MULTS_4_4(38)(PERCISION) & MULTS_4_4(38)(PERCISION downto 1));
			MULTS_5_2(39)<=signed(MULTS_4_3(39)(PERCISION) & MULTS_4_3(39)(PERCISION downto 1))+signed(MULTS_4_4(39)(PERCISION) & MULTS_4_4(39)(PERCISION downto 1));
			MULTS_5_2(40)<=signed(MULTS_4_3(40)(PERCISION) & MULTS_4_3(40)(PERCISION downto 1))+signed(MULTS_4_4(40)(PERCISION) & MULTS_4_4(40)(PERCISION downto 1));
			MULTS_5_2(41)<=signed(MULTS_4_3(41)(PERCISION) & MULTS_4_3(41)(PERCISION downto 1))+signed(MULTS_4_4(41)(PERCISION) & MULTS_4_4(41)(PERCISION downto 1));
			MULTS_5_2(42)<=signed(MULTS_4_3(42)(PERCISION) & MULTS_4_3(42)(PERCISION downto 1))+signed(MULTS_4_4(42)(PERCISION) & MULTS_4_4(42)(PERCISION downto 1));
			MULTS_5_2(43)<=signed(MULTS_4_3(43)(PERCISION) & MULTS_4_3(43)(PERCISION downto 1))+signed(MULTS_4_4(43)(PERCISION) & MULTS_4_4(43)(PERCISION downto 1));
			MULTS_5_2(44)<=signed(MULTS_4_3(44)(PERCISION) & MULTS_4_3(44)(PERCISION downto 1))+signed(MULTS_4_4(44)(PERCISION) & MULTS_4_4(44)(PERCISION downto 1));
			MULTS_5_2(45)<=signed(MULTS_4_3(45)(PERCISION) & MULTS_4_3(45)(PERCISION downto 1))+signed(MULTS_4_4(45)(PERCISION) & MULTS_4_4(45)(PERCISION downto 1));
			MULTS_5_2(46)<=signed(MULTS_4_3(46)(PERCISION) & MULTS_4_3(46)(PERCISION downto 1))+signed(MULTS_4_4(46)(PERCISION) & MULTS_4_4(46)(PERCISION downto 1));
			MULTS_5_2(47)<=signed(MULTS_4_3(47)(PERCISION) & MULTS_4_3(47)(PERCISION downto 1))+signed(MULTS_4_4(47)(PERCISION) & MULTS_4_4(47)(PERCISION downto 1));
			MULTS_5_2(48)<=signed(MULTS_4_3(48)(PERCISION) & MULTS_4_3(48)(PERCISION downto 1))+signed(MULTS_4_4(48)(PERCISION) & MULTS_4_4(48)(PERCISION downto 1));
			MULTS_5_2(49)<=signed(MULTS_4_3(49)(PERCISION) & MULTS_4_3(49)(PERCISION downto 1))+signed(MULTS_4_4(49)(PERCISION) & MULTS_4_4(49)(PERCISION downto 1));
			MULTS_5_2(50)<=signed(MULTS_4_3(50)(PERCISION) & MULTS_4_3(50)(PERCISION downto 1))+signed(MULTS_4_4(50)(PERCISION) & MULTS_4_4(50)(PERCISION downto 1));
			MULTS_5_2(51)<=signed(MULTS_4_3(51)(PERCISION) & MULTS_4_3(51)(PERCISION downto 1))+signed(MULTS_4_4(51)(PERCISION) & MULTS_4_4(51)(PERCISION downto 1));
			MULTS_5_2(52)<=signed(MULTS_4_3(52)(PERCISION) & MULTS_4_3(52)(PERCISION downto 1))+signed(MULTS_4_4(52)(PERCISION) & MULTS_4_4(52)(PERCISION downto 1));
			MULTS_5_2(53)<=signed(MULTS_4_3(53)(PERCISION) & MULTS_4_3(53)(PERCISION downto 1))+signed(MULTS_4_4(53)(PERCISION) & MULTS_4_4(53)(PERCISION downto 1));
			MULTS_5_2(54)<=signed(MULTS_4_3(54)(PERCISION) & MULTS_4_3(54)(PERCISION downto 1))+signed(MULTS_4_4(54)(PERCISION) & MULTS_4_4(54)(PERCISION downto 1));
			MULTS_5_2(55)<=signed(MULTS_4_3(55)(PERCISION) & MULTS_4_3(55)(PERCISION downto 1))+signed(MULTS_4_4(55)(PERCISION) & MULTS_4_4(55)(PERCISION downto 1));
			MULTS_5_2(56)<=signed(MULTS_4_3(56)(PERCISION) & MULTS_4_3(56)(PERCISION downto 1))+signed(MULTS_4_4(56)(PERCISION) & MULTS_4_4(56)(PERCISION downto 1));
			MULTS_5_2(57)<=signed(MULTS_4_3(57)(PERCISION) & MULTS_4_3(57)(PERCISION downto 1))+signed(MULTS_4_4(57)(PERCISION) & MULTS_4_4(57)(PERCISION downto 1));
			MULTS_5_2(58)<=signed(MULTS_4_3(58)(PERCISION) & MULTS_4_3(58)(PERCISION downto 1))+signed(MULTS_4_4(58)(PERCISION) & MULTS_4_4(58)(PERCISION downto 1));
			MULTS_5_2(59)<=signed(MULTS_4_3(59)(PERCISION) & MULTS_4_3(59)(PERCISION downto 1))+signed(MULTS_4_4(59)(PERCISION) & MULTS_4_4(59)(PERCISION downto 1));
			MULTS_5_2(60)<=signed(MULTS_4_3(60)(PERCISION) & MULTS_4_3(60)(PERCISION downto 1))+signed(MULTS_4_4(60)(PERCISION) & MULTS_4_4(60)(PERCISION downto 1));
			MULTS_5_2(61)<=signed(MULTS_4_3(61)(PERCISION) & MULTS_4_3(61)(PERCISION downto 1))+signed(MULTS_4_4(61)(PERCISION) & MULTS_4_4(61)(PERCISION downto 1));
			MULTS_5_2(62)<=signed(MULTS_4_3(62)(PERCISION) & MULTS_4_3(62)(PERCISION downto 1))+signed(MULTS_4_4(62)(PERCISION) & MULTS_4_4(62)(PERCISION downto 1));
			MULTS_5_2(63)<=signed(MULTS_4_3(63)(PERCISION) & MULTS_4_3(63)(PERCISION downto 1))+signed(MULTS_4_4(63)(PERCISION) & MULTS_4_4(63)(PERCISION downto 1));
			MULTS_5_2(64)<=signed(MULTS_4_3(64)(PERCISION) & MULTS_4_3(64)(PERCISION downto 1))+signed(MULTS_4_4(64)(PERCISION) & MULTS_4_4(64)(PERCISION downto 1));
			MULTS_5_2(65)<=signed(MULTS_4_3(65)(PERCISION) & MULTS_4_3(65)(PERCISION downto 1))+signed(MULTS_4_4(65)(PERCISION) & MULTS_4_4(65)(PERCISION downto 1));
			MULTS_5_2(66)<=signed(MULTS_4_3(66)(PERCISION) & MULTS_4_3(66)(PERCISION downto 1))+signed(MULTS_4_4(66)(PERCISION) & MULTS_4_4(66)(PERCISION downto 1));
			MULTS_5_2(67)<=signed(MULTS_4_3(67)(PERCISION) & MULTS_4_3(67)(PERCISION downto 1))+signed(MULTS_4_4(67)(PERCISION) & MULTS_4_4(67)(PERCISION downto 1));
			MULTS_5_2(68)<=signed(MULTS_4_3(68)(PERCISION) & MULTS_4_3(68)(PERCISION downto 1))+signed(MULTS_4_4(68)(PERCISION) & MULTS_4_4(68)(PERCISION downto 1));
			MULTS_5_2(69)<=signed(MULTS_4_3(69)(PERCISION) & MULTS_4_3(69)(PERCISION downto 1))+signed(MULTS_4_4(69)(PERCISION) & MULTS_4_4(69)(PERCISION downto 1));
			MULTS_5_2(70)<=signed(MULTS_4_3(70)(PERCISION) & MULTS_4_3(70)(PERCISION downto 1))+signed(MULTS_4_4(70)(PERCISION) & MULTS_4_4(70)(PERCISION downto 1));
			MULTS_5_2(71)<=signed(MULTS_4_3(71)(PERCISION) & MULTS_4_3(71)(PERCISION downto 1))+signed(MULTS_4_4(71)(PERCISION) & MULTS_4_4(71)(PERCISION downto 1));
			MULTS_5_2(72)<=signed(MULTS_4_3(72)(PERCISION) & MULTS_4_3(72)(PERCISION downto 1))+signed(MULTS_4_4(72)(PERCISION) & MULTS_4_4(72)(PERCISION downto 1));
			MULTS_5_2(73)<=signed(MULTS_4_3(73)(PERCISION) & MULTS_4_3(73)(PERCISION downto 1))+signed(MULTS_4_4(73)(PERCISION) & MULTS_4_4(73)(PERCISION downto 1));
			MULTS_5_2(74)<=signed(MULTS_4_3(74)(PERCISION) & MULTS_4_3(74)(PERCISION downto 1))+signed(MULTS_4_4(74)(PERCISION) & MULTS_4_4(74)(PERCISION downto 1));
			MULTS_5_2(75)<=signed(MULTS_4_3(75)(PERCISION) & MULTS_4_3(75)(PERCISION downto 1))+signed(MULTS_4_4(75)(PERCISION) & MULTS_4_4(75)(PERCISION downto 1));
			MULTS_5_2(76)<=signed(MULTS_4_3(76)(PERCISION) & MULTS_4_3(76)(PERCISION downto 1))+signed(MULTS_4_4(76)(PERCISION) & MULTS_4_4(76)(PERCISION downto 1));
			MULTS_5_2(77)<=signed(MULTS_4_3(77)(PERCISION) & MULTS_4_3(77)(PERCISION downto 1))+signed(MULTS_4_4(77)(PERCISION) & MULTS_4_4(77)(PERCISION downto 1));
			MULTS_5_2(78)<=signed(MULTS_4_3(78)(PERCISION) & MULTS_4_3(78)(PERCISION downto 1))+signed(MULTS_4_4(78)(PERCISION) & MULTS_4_4(78)(PERCISION downto 1));
			MULTS_5_2(79)<=signed(MULTS_4_3(79)(PERCISION) & MULTS_4_3(79)(PERCISION downto 1))+signed(MULTS_4_4(79)(PERCISION) & MULTS_4_4(79)(PERCISION downto 1));
			MULTS_5_2(80)<=signed(MULTS_4_3(80)(PERCISION) & MULTS_4_3(80)(PERCISION downto 1))+signed(MULTS_4_4(80)(PERCISION) & MULTS_4_4(80)(PERCISION downto 1));
			MULTS_5_2(81)<=signed(MULTS_4_3(81)(PERCISION) & MULTS_4_3(81)(PERCISION downto 1))+signed(MULTS_4_4(81)(PERCISION) & MULTS_4_4(81)(PERCISION downto 1));
			MULTS_5_2(82)<=signed(MULTS_4_3(82)(PERCISION) & MULTS_4_3(82)(PERCISION downto 1))+signed(MULTS_4_4(82)(PERCISION) & MULTS_4_4(82)(PERCISION downto 1));
			MULTS_5_2(83)<=signed(MULTS_4_3(83)(PERCISION) & MULTS_4_3(83)(PERCISION downto 1))+signed(MULTS_4_4(83)(PERCISION) & MULTS_4_4(83)(PERCISION downto 1));



                         EN_SUM_MULT_6<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_6 = '1' then
			------------------------------------STAGE-6--------------------------------------
			MULTS_6_1(0)<=signed(MULTS_5_1(0)(PERCISION) & MULTS_5_1(0)(PERCISION downto 1))+signed(MULTS_5_2(0)(PERCISION) & MULTS_5_2(0)(PERCISION downto 1));
			MULTS_6_1(1)<=signed(MULTS_5_1(1)(PERCISION) & MULTS_5_1(1)(PERCISION downto 1))+signed(MULTS_5_2(1)(PERCISION) & MULTS_5_2(1)(PERCISION downto 1));
			MULTS_6_1(2)<=signed(MULTS_5_1(2)(PERCISION) & MULTS_5_1(2)(PERCISION downto 1))+signed(MULTS_5_2(2)(PERCISION) & MULTS_5_2(2)(PERCISION downto 1));
			MULTS_6_1(3)<=signed(MULTS_5_1(3)(PERCISION) & MULTS_5_1(3)(PERCISION downto 1))+signed(MULTS_5_2(3)(PERCISION) & MULTS_5_2(3)(PERCISION downto 1));
			MULTS_6_1(4)<=signed(MULTS_5_1(4)(PERCISION) & MULTS_5_1(4)(PERCISION downto 1))+signed(MULTS_5_2(4)(PERCISION) & MULTS_5_2(4)(PERCISION downto 1));
			MULTS_6_1(5)<=signed(MULTS_5_1(5)(PERCISION) & MULTS_5_1(5)(PERCISION downto 1))+signed(MULTS_5_2(5)(PERCISION) & MULTS_5_2(5)(PERCISION downto 1));
			MULTS_6_1(6)<=signed(MULTS_5_1(6)(PERCISION) & MULTS_5_1(6)(PERCISION downto 1))+signed(MULTS_5_2(6)(PERCISION) & MULTS_5_2(6)(PERCISION downto 1));
			MULTS_6_1(7)<=signed(MULTS_5_1(7)(PERCISION) & MULTS_5_1(7)(PERCISION downto 1))+signed(MULTS_5_2(7)(PERCISION) & MULTS_5_2(7)(PERCISION downto 1));
			MULTS_6_1(8)<=signed(MULTS_5_1(8)(PERCISION) & MULTS_5_1(8)(PERCISION downto 1))+signed(MULTS_5_2(8)(PERCISION) & MULTS_5_2(8)(PERCISION downto 1));
			MULTS_6_1(9)<=signed(MULTS_5_1(9)(PERCISION) & MULTS_5_1(9)(PERCISION downto 1))+signed(MULTS_5_2(9)(PERCISION) & MULTS_5_2(9)(PERCISION downto 1));
			MULTS_6_1(10)<=signed(MULTS_5_1(10)(PERCISION) & MULTS_5_1(10)(PERCISION downto 1))+signed(MULTS_5_2(10)(PERCISION) & MULTS_5_2(10)(PERCISION downto 1));
			MULTS_6_1(11)<=signed(MULTS_5_1(11)(PERCISION) & MULTS_5_1(11)(PERCISION downto 1))+signed(MULTS_5_2(11)(PERCISION) & MULTS_5_2(11)(PERCISION downto 1));
			MULTS_6_1(12)<=signed(MULTS_5_1(12)(PERCISION) & MULTS_5_1(12)(PERCISION downto 1))+signed(MULTS_5_2(12)(PERCISION) & MULTS_5_2(12)(PERCISION downto 1));
			MULTS_6_1(13)<=signed(MULTS_5_1(13)(PERCISION) & MULTS_5_1(13)(PERCISION downto 1))+signed(MULTS_5_2(13)(PERCISION) & MULTS_5_2(13)(PERCISION downto 1));
			MULTS_6_1(14)<=signed(MULTS_5_1(14)(PERCISION) & MULTS_5_1(14)(PERCISION downto 1))+signed(MULTS_5_2(14)(PERCISION) & MULTS_5_2(14)(PERCISION downto 1));
			MULTS_6_1(15)<=signed(MULTS_5_1(15)(PERCISION) & MULTS_5_1(15)(PERCISION downto 1))+signed(MULTS_5_2(15)(PERCISION) & MULTS_5_2(15)(PERCISION downto 1));
			MULTS_6_1(16)<=signed(MULTS_5_1(16)(PERCISION) & MULTS_5_1(16)(PERCISION downto 1))+signed(MULTS_5_2(16)(PERCISION) & MULTS_5_2(16)(PERCISION downto 1));
			MULTS_6_1(17)<=signed(MULTS_5_1(17)(PERCISION) & MULTS_5_1(17)(PERCISION downto 1))+signed(MULTS_5_2(17)(PERCISION) & MULTS_5_2(17)(PERCISION downto 1));
			MULTS_6_1(18)<=signed(MULTS_5_1(18)(PERCISION) & MULTS_5_1(18)(PERCISION downto 1))+signed(MULTS_5_2(18)(PERCISION) & MULTS_5_2(18)(PERCISION downto 1));
			MULTS_6_1(19)<=signed(MULTS_5_1(19)(PERCISION) & MULTS_5_1(19)(PERCISION downto 1))+signed(MULTS_5_2(19)(PERCISION) & MULTS_5_2(19)(PERCISION downto 1));
			MULTS_6_1(20)<=signed(MULTS_5_1(20)(PERCISION) & MULTS_5_1(20)(PERCISION downto 1))+signed(MULTS_5_2(20)(PERCISION) & MULTS_5_2(20)(PERCISION downto 1));
			MULTS_6_1(21)<=signed(MULTS_5_1(21)(PERCISION) & MULTS_5_1(21)(PERCISION downto 1))+signed(MULTS_5_2(21)(PERCISION) & MULTS_5_2(21)(PERCISION downto 1));
			MULTS_6_1(22)<=signed(MULTS_5_1(22)(PERCISION) & MULTS_5_1(22)(PERCISION downto 1))+signed(MULTS_5_2(22)(PERCISION) & MULTS_5_2(22)(PERCISION downto 1));
			MULTS_6_1(23)<=signed(MULTS_5_1(23)(PERCISION) & MULTS_5_1(23)(PERCISION downto 1))+signed(MULTS_5_2(23)(PERCISION) & MULTS_5_2(23)(PERCISION downto 1));
			MULTS_6_1(24)<=signed(MULTS_5_1(24)(PERCISION) & MULTS_5_1(24)(PERCISION downto 1))+signed(MULTS_5_2(24)(PERCISION) & MULTS_5_2(24)(PERCISION downto 1));
			MULTS_6_1(25)<=signed(MULTS_5_1(25)(PERCISION) & MULTS_5_1(25)(PERCISION downto 1))+signed(MULTS_5_2(25)(PERCISION) & MULTS_5_2(25)(PERCISION downto 1));
			MULTS_6_1(26)<=signed(MULTS_5_1(26)(PERCISION) & MULTS_5_1(26)(PERCISION downto 1))+signed(MULTS_5_2(26)(PERCISION) & MULTS_5_2(26)(PERCISION downto 1));
			MULTS_6_1(27)<=signed(MULTS_5_1(27)(PERCISION) & MULTS_5_1(27)(PERCISION downto 1))+signed(MULTS_5_2(27)(PERCISION) & MULTS_5_2(27)(PERCISION downto 1));
			MULTS_6_1(28)<=signed(MULTS_5_1(28)(PERCISION) & MULTS_5_1(28)(PERCISION downto 1))+signed(MULTS_5_2(28)(PERCISION) & MULTS_5_2(28)(PERCISION downto 1));
			MULTS_6_1(29)<=signed(MULTS_5_1(29)(PERCISION) & MULTS_5_1(29)(PERCISION downto 1))+signed(MULTS_5_2(29)(PERCISION) & MULTS_5_2(29)(PERCISION downto 1));
			MULTS_6_1(30)<=signed(MULTS_5_1(30)(PERCISION) & MULTS_5_1(30)(PERCISION downto 1))+signed(MULTS_5_2(30)(PERCISION) & MULTS_5_2(30)(PERCISION downto 1));
			MULTS_6_1(31)<=signed(MULTS_5_1(31)(PERCISION) & MULTS_5_1(31)(PERCISION downto 1))+signed(MULTS_5_2(31)(PERCISION) & MULTS_5_2(31)(PERCISION downto 1));
			MULTS_6_1(32)<=signed(MULTS_5_1(32)(PERCISION) & MULTS_5_1(32)(PERCISION downto 1))+signed(MULTS_5_2(32)(PERCISION) & MULTS_5_2(32)(PERCISION downto 1));
			MULTS_6_1(33)<=signed(MULTS_5_1(33)(PERCISION) & MULTS_5_1(33)(PERCISION downto 1))+signed(MULTS_5_2(33)(PERCISION) & MULTS_5_2(33)(PERCISION downto 1));
			MULTS_6_1(34)<=signed(MULTS_5_1(34)(PERCISION) & MULTS_5_1(34)(PERCISION downto 1))+signed(MULTS_5_2(34)(PERCISION) & MULTS_5_2(34)(PERCISION downto 1));
			MULTS_6_1(35)<=signed(MULTS_5_1(35)(PERCISION) & MULTS_5_1(35)(PERCISION downto 1))+signed(MULTS_5_2(35)(PERCISION) & MULTS_5_2(35)(PERCISION downto 1));
			MULTS_6_1(36)<=signed(MULTS_5_1(36)(PERCISION) & MULTS_5_1(36)(PERCISION downto 1))+signed(MULTS_5_2(36)(PERCISION) & MULTS_5_2(36)(PERCISION downto 1));
			MULTS_6_1(37)<=signed(MULTS_5_1(37)(PERCISION) & MULTS_5_1(37)(PERCISION downto 1))+signed(MULTS_5_2(37)(PERCISION) & MULTS_5_2(37)(PERCISION downto 1));
			MULTS_6_1(38)<=signed(MULTS_5_1(38)(PERCISION) & MULTS_5_1(38)(PERCISION downto 1))+signed(MULTS_5_2(38)(PERCISION) & MULTS_5_2(38)(PERCISION downto 1));
			MULTS_6_1(39)<=signed(MULTS_5_1(39)(PERCISION) & MULTS_5_1(39)(PERCISION downto 1))+signed(MULTS_5_2(39)(PERCISION) & MULTS_5_2(39)(PERCISION downto 1));
			MULTS_6_1(40)<=signed(MULTS_5_1(40)(PERCISION) & MULTS_5_1(40)(PERCISION downto 1))+signed(MULTS_5_2(40)(PERCISION) & MULTS_5_2(40)(PERCISION downto 1));
			MULTS_6_1(41)<=signed(MULTS_5_1(41)(PERCISION) & MULTS_5_1(41)(PERCISION downto 1))+signed(MULTS_5_2(41)(PERCISION) & MULTS_5_2(41)(PERCISION downto 1));
			MULTS_6_1(42)<=signed(MULTS_5_1(42)(PERCISION) & MULTS_5_1(42)(PERCISION downto 1))+signed(MULTS_5_2(42)(PERCISION) & MULTS_5_2(42)(PERCISION downto 1));
			MULTS_6_1(43)<=signed(MULTS_5_1(43)(PERCISION) & MULTS_5_1(43)(PERCISION downto 1))+signed(MULTS_5_2(43)(PERCISION) & MULTS_5_2(43)(PERCISION downto 1));
			MULTS_6_1(44)<=signed(MULTS_5_1(44)(PERCISION) & MULTS_5_1(44)(PERCISION downto 1))+signed(MULTS_5_2(44)(PERCISION) & MULTS_5_2(44)(PERCISION downto 1));
			MULTS_6_1(45)<=signed(MULTS_5_1(45)(PERCISION) & MULTS_5_1(45)(PERCISION downto 1))+signed(MULTS_5_2(45)(PERCISION) & MULTS_5_2(45)(PERCISION downto 1));
			MULTS_6_1(46)<=signed(MULTS_5_1(46)(PERCISION) & MULTS_5_1(46)(PERCISION downto 1))+signed(MULTS_5_2(46)(PERCISION) & MULTS_5_2(46)(PERCISION downto 1));
			MULTS_6_1(47)<=signed(MULTS_5_1(47)(PERCISION) & MULTS_5_1(47)(PERCISION downto 1))+signed(MULTS_5_2(47)(PERCISION) & MULTS_5_2(47)(PERCISION downto 1));
			MULTS_6_1(48)<=signed(MULTS_5_1(48)(PERCISION) & MULTS_5_1(48)(PERCISION downto 1))+signed(MULTS_5_2(48)(PERCISION) & MULTS_5_2(48)(PERCISION downto 1));
			MULTS_6_1(49)<=signed(MULTS_5_1(49)(PERCISION) & MULTS_5_1(49)(PERCISION downto 1))+signed(MULTS_5_2(49)(PERCISION) & MULTS_5_2(49)(PERCISION downto 1));
			MULTS_6_1(50)<=signed(MULTS_5_1(50)(PERCISION) & MULTS_5_1(50)(PERCISION downto 1))+signed(MULTS_5_2(50)(PERCISION) & MULTS_5_2(50)(PERCISION downto 1));
			MULTS_6_1(51)<=signed(MULTS_5_1(51)(PERCISION) & MULTS_5_1(51)(PERCISION downto 1))+signed(MULTS_5_2(51)(PERCISION) & MULTS_5_2(51)(PERCISION downto 1));
			MULTS_6_1(52)<=signed(MULTS_5_1(52)(PERCISION) & MULTS_5_1(52)(PERCISION downto 1))+signed(MULTS_5_2(52)(PERCISION) & MULTS_5_2(52)(PERCISION downto 1));
			MULTS_6_1(53)<=signed(MULTS_5_1(53)(PERCISION) & MULTS_5_1(53)(PERCISION downto 1))+signed(MULTS_5_2(53)(PERCISION) & MULTS_5_2(53)(PERCISION downto 1));
			MULTS_6_1(54)<=signed(MULTS_5_1(54)(PERCISION) & MULTS_5_1(54)(PERCISION downto 1))+signed(MULTS_5_2(54)(PERCISION) & MULTS_5_2(54)(PERCISION downto 1));
			MULTS_6_1(55)<=signed(MULTS_5_1(55)(PERCISION) & MULTS_5_1(55)(PERCISION downto 1))+signed(MULTS_5_2(55)(PERCISION) & MULTS_5_2(55)(PERCISION downto 1));
			MULTS_6_1(56)<=signed(MULTS_5_1(56)(PERCISION) & MULTS_5_1(56)(PERCISION downto 1))+signed(MULTS_5_2(56)(PERCISION) & MULTS_5_2(56)(PERCISION downto 1));
			MULTS_6_1(57)<=signed(MULTS_5_1(57)(PERCISION) & MULTS_5_1(57)(PERCISION downto 1))+signed(MULTS_5_2(57)(PERCISION) & MULTS_5_2(57)(PERCISION downto 1));
			MULTS_6_1(58)<=signed(MULTS_5_1(58)(PERCISION) & MULTS_5_1(58)(PERCISION downto 1))+signed(MULTS_5_2(58)(PERCISION) & MULTS_5_2(58)(PERCISION downto 1));
			MULTS_6_1(59)<=signed(MULTS_5_1(59)(PERCISION) & MULTS_5_1(59)(PERCISION downto 1))+signed(MULTS_5_2(59)(PERCISION) & MULTS_5_2(59)(PERCISION downto 1));
			MULTS_6_1(60)<=signed(MULTS_5_1(60)(PERCISION) & MULTS_5_1(60)(PERCISION downto 1))+signed(MULTS_5_2(60)(PERCISION) & MULTS_5_2(60)(PERCISION downto 1));
			MULTS_6_1(61)<=signed(MULTS_5_1(61)(PERCISION) & MULTS_5_1(61)(PERCISION downto 1))+signed(MULTS_5_2(61)(PERCISION) & MULTS_5_2(61)(PERCISION downto 1));
			MULTS_6_1(62)<=signed(MULTS_5_1(62)(PERCISION) & MULTS_5_1(62)(PERCISION downto 1))+signed(MULTS_5_2(62)(PERCISION) & MULTS_5_2(62)(PERCISION downto 1));
			MULTS_6_1(63)<=signed(MULTS_5_1(63)(PERCISION) & MULTS_5_1(63)(PERCISION downto 1))+signed(MULTS_5_2(63)(PERCISION) & MULTS_5_2(63)(PERCISION downto 1));
			MULTS_6_1(64)<=signed(MULTS_5_1(64)(PERCISION) & MULTS_5_1(64)(PERCISION downto 1))+signed(MULTS_5_2(64)(PERCISION) & MULTS_5_2(64)(PERCISION downto 1));
			MULTS_6_1(65)<=signed(MULTS_5_1(65)(PERCISION) & MULTS_5_1(65)(PERCISION downto 1))+signed(MULTS_5_2(65)(PERCISION) & MULTS_5_2(65)(PERCISION downto 1));
			MULTS_6_1(66)<=signed(MULTS_5_1(66)(PERCISION) & MULTS_5_1(66)(PERCISION downto 1))+signed(MULTS_5_2(66)(PERCISION) & MULTS_5_2(66)(PERCISION downto 1));
			MULTS_6_1(67)<=signed(MULTS_5_1(67)(PERCISION) & MULTS_5_1(67)(PERCISION downto 1))+signed(MULTS_5_2(67)(PERCISION) & MULTS_5_2(67)(PERCISION downto 1));
			MULTS_6_1(68)<=signed(MULTS_5_1(68)(PERCISION) & MULTS_5_1(68)(PERCISION downto 1))+signed(MULTS_5_2(68)(PERCISION) & MULTS_5_2(68)(PERCISION downto 1));
			MULTS_6_1(69)<=signed(MULTS_5_1(69)(PERCISION) & MULTS_5_1(69)(PERCISION downto 1))+signed(MULTS_5_2(69)(PERCISION) & MULTS_5_2(69)(PERCISION downto 1));
			MULTS_6_1(70)<=signed(MULTS_5_1(70)(PERCISION) & MULTS_5_1(70)(PERCISION downto 1))+signed(MULTS_5_2(70)(PERCISION) & MULTS_5_2(70)(PERCISION downto 1));
			MULTS_6_1(71)<=signed(MULTS_5_1(71)(PERCISION) & MULTS_5_1(71)(PERCISION downto 1))+signed(MULTS_5_2(71)(PERCISION) & MULTS_5_2(71)(PERCISION downto 1));
			MULTS_6_1(72)<=signed(MULTS_5_1(72)(PERCISION) & MULTS_5_1(72)(PERCISION downto 1))+signed(MULTS_5_2(72)(PERCISION) & MULTS_5_2(72)(PERCISION downto 1));
			MULTS_6_1(73)<=signed(MULTS_5_1(73)(PERCISION) & MULTS_5_1(73)(PERCISION downto 1))+signed(MULTS_5_2(73)(PERCISION) & MULTS_5_2(73)(PERCISION downto 1));
			MULTS_6_1(74)<=signed(MULTS_5_1(74)(PERCISION) & MULTS_5_1(74)(PERCISION downto 1))+signed(MULTS_5_2(74)(PERCISION) & MULTS_5_2(74)(PERCISION downto 1));
			MULTS_6_1(75)<=signed(MULTS_5_1(75)(PERCISION) & MULTS_5_1(75)(PERCISION downto 1))+signed(MULTS_5_2(75)(PERCISION) & MULTS_5_2(75)(PERCISION downto 1));
			MULTS_6_1(76)<=signed(MULTS_5_1(76)(PERCISION) & MULTS_5_1(76)(PERCISION downto 1))+signed(MULTS_5_2(76)(PERCISION) & MULTS_5_2(76)(PERCISION downto 1));
			MULTS_6_1(77)<=signed(MULTS_5_1(77)(PERCISION) & MULTS_5_1(77)(PERCISION downto 1))+signed(MULTS_5_2(77)(PERCISION) & MULTS_5_2(77)(PERCISION downto 1));
			MULTS_6_1(78)<=signed(MULTS_5_1(78)(PERCISION) & MULTS_5_1(78)(PERCISION downto 1))+signed(MULTS_5_2(78)(PERCISION) & MULTS_5_2(78)(PERCISION downto 1));
			MULTS_6_1(79)<=signed(MULTS_5_1(79)(PERCISION) & MULTS_5_1(79)(PERCISION downto 1))+signed(MULTS_5_2(79)(PERCISION) & MULTS_5_2(79)(PERCISION downto 1));
			MULTS_6_1(80)<=signed(MULTS_5_1(80)(PERCISION) & MULTS_5_1(80)(PERCISION downto 1))+signed(MULTS_5_2(80)(PERCISION) & MULTS_5_2(80)(PERCISION downto 1));
			MULTS_6_1(81)<=signed(MULTS_5_1(81)(PERCISION) & MULTS_5_1(81)(PERCISION downto 1))+signed(MULTS_5_2(81)(PERCISION) & MULTS_5_2(81)(PERCISION downto 1));
			MULTS_6_1(82)<=signed(MULTS_5_1(82)(PERCISION) & MULTS_5_1(82)(PERCISION downto 1))+signed(MULTS_5_2(82)(PERCISION) & MULTS_5_2(82)(PERCISION downto 1));
			MULTS_6_1(83)<=signed(MULTS_5_1(83)(PERCISION) & MULTS_5_1(83)(PERCISION downto 1))+signed(MULTS_5_2(83)(PERCISION) & MULTS_5_2(83)(PERCISION downto 1));



                         EN_SUM_MULT_7<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_7 = '1' then
			------------------------------------STAGE-7--------------------------------------
			MULTS_7_1(0)<=signed(MULTS_6_1(0)(PERCISION) & MULTS_6_1(0)(PERCISION downto 1))+signed(MULTS_6_2(0)(PERCISION) & MULTS_6_2(0)(PERCISION downto 1));
			MULTS_7_1(1)<=signed(MULTS_6_1(1)(PERCISION) & MULTS_6_1(1)(PERCISION downto 1))+signed(MULTS_6_2(1)(PERCISION) & MULTS_6_2(1)(PERCISION downto 1));
			MULTS_7_1(2)<=signed(MULTS_6_1(2)(PERCISION) & MULTS_6_1(2)(PERCISION downto 1))+signed(MULTS_6_2(2)(PERCISION) & MULTS_6_2(2)(PERCISION downto 1));
			MULTS_7_1(3)<=signed(MULTS_6_1(3)(PERCISION) & MULTS_6_1(3)(PERCISION downto 1))+signed(MULTS_6_2(3)(PERCISION) & MULTS_6_2(3)(PERCISION downto 1));
			MULTS_7_1(4)<=signed(MULTS_6_1(4)(PERCISION) & MULTS_6_1(4)(PERCISION downto 1))+signed(MULTS_6_2(4)(PERCISION) & MULTS_6_2(4)(PERCISION downto 1));
			MULTS_7_1(5)<=signed(MULTS_6_1(5)(PERCISION) & MULTS_6_1(5)(PERCISION downto 1))+signed(MULTS_6_2(5)(PERCISION) & MULTS_6_2(5)(PERCISION downto 1));
			MULTS_7_1(6)<=signed(MULTS_6_1(6)(PERCISION) & MULTS_6_1(6)(PERCISION downto 1))+signed(MULTS_6_2(6)(PERCISION) & MULTS_6_2(6)(PERCISION downto 1));
			MULTS_7_1(7)<=signed(MULTS_6_1(7)(PERCISION) & MULTS_6_1(7)(PERCISION downto 1))+signed(MULTS_6_2(7)(PERCISION) & MULTS_6_2(7)(PERCISION downto 1));
			MULTS_7_1(8)<=signed(MULTS_6_1(8)(PERCISION) & MULTS_6_1(8)(PERCISION downto 1))+signed(MULTS_6_2(8)(PERCISION) & MULTS_6_2(8)(PERCISION downto 1));
			MULTS_7_1(9)<=signed(MULTS_6_1(9)(PERCISION) & MULTS_6_1(9)(PERCISION downto 1))+signed(MULTS_6_2(9)(PERCISION) & MULTS_6_2(9)(PERCISION downto 1));
			MULTS_7_1(10)<=signed(MULTS_6_1(10)(PERCISION) & MULTS_6_1(10)(PERCISION downto 1))+signed(MULTS_6_2(10)(PERCISION) & MULTS_6_2(10)(PERCISION downto 1));
			MULTS_7_1(11)<=signed(MULTS_6_1(11)(PERCISION) & MULTS_6_1(11)(PERCISION downto 1))+signed(MULTS_6_2(11)(PERCISION) & MULTS_6_2(11)(PERCISION downto 1));
			MULTS_7_1(12)<=signed(MULTS_6_1(12)(PERCISION) & MULTS_6_1(12)(PERCISION downto 1))+signed(MULTS_6_2(12)(PERCISION) & MULTS_6_2(12)(PERCISION downto 1));
			MULTS_7_1(13)<=signed(MULTS_6_1(13)(PERCISION) & MULTS_6_1(13)(PERCISION downto 1))+signed(MULTS_6_2(13)(PERCISION) & MULTS_6_2(13)(PERCISION downto 1));
			MULTS_7_1(14)<=signed(MULTS_6_1(14)(PERCISION) & MULTS_6_1(14)(PERCISION downto 1))+signed(MULTS_6_2(14)(PERCISION) & MULTS_6_2(14)(PERCISION downto 1));
			MULTS_7_1(15)<=signed(MULTS_6_1(15)(PERCISION) & MULTS_6_1(15)(PERCISION downto 1))+signed(MULTS_6_2(15)(PERCISION) & MULTS_6_2(15)(PERCISION downto 1));
			MULTS_7_1(16)<=signed(MULTS_6_1(16)(PERCISION) & MULTS_6_1(16)(PERCISION downto 1))+signed(MULTS_6_2(16)(PERCISION) & MULTS_6_2(16)(PERCISION downto 1));
			MULTS_7_1(17)<=signed(MULTS_6_1(17)(PERCISION) & MULTS_6_1(17)(PERCISION downto 1))+signed(MULTS_6_2(17)(PERCISION) & MULTS_6_2(17)(PERCISION downto 1));
			MULTS_7_1(18)<=signed(MULTS_6_1(18)(PERCISION) & MULTS_6_1(18)(PERCISION downto 1))+signed(MULTS_6_2(18)(PERCISION) & MULTS_6_2(18)(PERCISION downto 1));
			MULTS_7_1(19)<=signed(MULTS_6_1(19)(PERCISION) & MULTS_6_1(19)(PERCISION downto 1))+signed(MULTS_6_2(19)(PERCISION) & MULTS_6_2(19)(PERCISION downto 1));
			MULTS_7_1(20)<=signed(MULTS_6_1(20)(PERCISION) & MULTS_6_1(20)(PERCISION downto 1))+signed(MULTS_6_2(20)(PERCISION) & MULTS_6_2(20)(PERCISION downto 1));
			MULTS_7_1(21)<=signed(MULTS_6_1(21)(PERCISION) & MULTS_6_1(21)(PERCISION downto 1))+signed(MULTS_6_2(21)(PERCISION) & MULTS_6_2(21)(PERCISION downto 1));
			MULTS_7_1(22)<=signed(MULTS_6_1(22)(PERCISION) & MULTS_6_1(22)(PERCISION downto 1))+signed(MULTS_6_2(22)(PERCISION) & MULTS_6_2(22)(PERCISION downto 1));
			MULTS_7_1(23)<=signed(MULTS_6_1(23)(PERCISION) & MULTS_6_1(23)(PERCISION downto 1))+signed(MULTS_6_2(23)(PERCISION) & MULTS_6_2(23)(PERCISION downto 1));
			MULTS_7_1(24)<=signed(MULTS_6_1(24)(PERCISION) & MULTS_6_1(24)(PERCISION downto 1))+signed(MULTS_6_2(24)(PERCISION) & MULTS_6_2(24)(PERCISION downto 1));
			MULTS_7_1(25)<=signed(MULTS_6_1(25)(PERCISION) & MULTS_6_1(25)(PERCISION downto 1))+signed(MULTS_6_2(25)(PERCISION) & MULTS_6_2(25)(PERCISION downto 1));
			MULTS_7_1(26)<=signed(MULTS_6_1(26)(PERCISION) & MULTS_6_1(26)(PERCISION downto 1))+signed(MULTS_6_2(26)(PERCISION) & MULTS_6_2(26)(PERCISION downto 1));
			MULTS_7_1(27)<=signed(MULTS_6_1(27)(PERCISION) & MULTS_6_1(27)(PERCISION downto 1))+signed(MULTS_6_2(27)(PERCISION) & MULTS_6_2(27)(PERCISION downto 1));
			MULTS_7_1(28)<=signed(MULTS_6_1(28)(PERCISION) & MULTS_6_1(28)(PERCISION downto 1))+signed(MULTS_6_2(28)(PERCISION) & MULTS_6_2(28)(PERCISION downto 1));
			MULTS_7_1(29)<=signed(MULTS_6_1(29)(PERCISION) & MULTS_6_1(29)(PERCISION downto 1))+signed(MULTS_6_2(29)(PERCISION) & MULTS_6_2(29)(PERCISION downto 1));
			MULTS_7_1(30)<=signed(MULTS_6_1(30)(PERCISION) & MULTS_6_1(30)(PERCISION downto 1))+signed(MULTS_6_2(30)(PERCISION) & MULTS_6_2(30)(PERCISION downto 1));
			MULTS_7_1(31)<=signed(MULTS_6_1(31)(PERCISION) & MULTS_6_1(31)(PERCISION downto 1))+signed(MULTS_6_2(31)(PERCISION) & MULTS_6_2(31)(PERCISION downto 1));
			MULTS_7_1(32)<=signed(MULTS_6_1(32)(PERCISION) & MULTS_6_1(32)(PERCISION downto 1))+signed(MULTS_6_2(32)(PERCISION) & MULTS_6_2(32)(PERCISION downto 1));
			MULTS_7_1(33)<=signed(MULTS_6_1(33)(PERCISION) & MULTS_6_1(33)(PERCISION downto 1))+signed(MULTS_6_2(33)(PERCISION) & MULTS_6_2(33)(PERCISION downto 1));
			MULTS_7_1(34)<=signed(MULTS_6_1(34)(PERCISION) & MULTS_6_1(34)(PERCISION downto 1))+signed(MULTS_6_2(34)(PERCISION) & MULTS_6_2(34)(PERCISION downto 1));
			MULTS_7_1(35)<=signed(MULTS_6_1(35)(PERCISION) & MULTS_6_1(35)(PERCISION downto 1))+signed(MULTS_6_2(35)(PERCISION) & MULTS_6_2(35)(PERCISION downto 1));
			MULTS_7_1(36)<=signed(MULTS_6_1(36)(PERCISION) & MULTS_6_1(36)(PERCISION downto 1))+signed(MULTS_6_2(36)(PERCISION) & MULTS_6_2(36)(PERCISION downto 1));
			MULTS_7_1(37)<=signed(MULTS_6_1(37)(PERCISION) & MULTS_6_1(37)(PERCISION downto 1))+signed(MULTS_6_2(37)(PERCISION) & MULTS_6_2(37)(PERCISION downto 1));
			MULTS_7_1(38)<=signed(MULTS_6_1(38)(PERCISION) & MULTS_6_1(38)(PERCISION downto 1))+signed(MULTS_6_2(38)(PERCISION) & MULTS_6_2(38)(PERCISION downto 1));
			MULTS_7_1(39)<=signed(MULTS_6_1(39)(PERCISION) & MULTS_6_1(39)(PERCISION downto 1))+signed(MULTS_6_2(39)(PERCISION) & MULTS_6_2(39)(PERCISION downto 1));
			MULTS_7_1(40)<=signed(MULTS_6_1(40)(PERCISION) & MULTS_6_1(40)(PERCISION downto 1))+signed(MULTS_6_2(40)(PERCISION) & MULTS_6_2(40)(PERCISION downto 1));
			MULTS_7_1(41)<=signed(MULTS_6_1(41)(PERCISION) & MULTS_6_1(41)(PERCISION downto 1))+signed(MULTS_6_2(41)(PERCISION) & MULTS_6_2(41)(PERCISION downto 1));
			MULTS_7_1(42)<=signed(MULTS_6_1(42)(PERCISION) & MULTS_6_1(42)(PERCISION downto 1))+signed(MULTS_6_2(42)(PERCISION) & MULTS_6_2(42)(PERCISION downto 1));
			MULTS_7_1(43)<=signed(MULTS_6_1(43)(PERCISION) & MULTS_6_1(43)(PERCISION downto 1))+signed(MULTS_6_2(43)(PERCISION) & MULTS_6_2(43)(PERCISION downto 1));
			MULTS_7_1(44)<=signed(MULTS_6_1(44)(PERCISION) & MULTS_6_1(44)(PERCISION downto 1))+signed(MULTS_6_2(44)(PERCISION) & MULTS_6_2(44)(PERCISION downto 1));
			MULTS_7_1(45)<=signed(MULTS_6_1(45)(PERCISION) & MULTS_6_1(45)(PERCISION downto 1))+signed(MULTS_6_2(45)(PERCISION) & MULTS_6_2(45)(PERCISION downto 1));
			MULTS_7_1(46)<=signed(MULTS_6_1(46)(PERCISION) & MULTS_6_1(46)(PERCISION downto 1))+signed(MULTS_6_2(46)(PERCISION) & MULTS_6_2(46)(PERCISION downto 1));
			MULTS_7_1(47)<=signed(MULTS_6_1(47)(PERCISION) & MULTS_6_1(47)(PERCISION downto 1))+signed(MULTS_6_2(47)(PERCISION) & MULTS_6_2(47)(PERCISION downto 1));
			MULTS_7_1(48)<=signed(MULTS_6_1(48)(PERCISION) & MULTS_6_1(48)(PERCISION downto 1))+signed(MULTS_6_2(48)(PERCISION) & MULTS_6_2(48)(PERCISION downto 1));
			MULTS_7_1(49)<=signed(MULTS_6_1(49)(PERCISION) & MULTS_6_1(49)(PERCISION downto 1))+signed(MULTS_6_2(49)(PERCISION) & MULTS_6_2(49)(PERCISION downto 1));
			MULTS_7_1(50)<=signed(MULTS_6_1(50)(PERCISION) & MULTS_6_1(50)(PERCISION downto 1))+signed(MULTS_6_2(50)(PERCISION) & MULTS_6_2(50)(PERCISION downto 1));
			MULTS_7_1(51)<=signed(MULTS_6_1(51)(PERCISION) & MULTS_6_1(51)(PERCISION downto 1))+signed(MULTS_6_2(51)(PERCISION) & MULTS_6_2(51)(PERCISION downto 1));
			MULTS_7_1(52)<=signed(MULTS_6_1(52)(PERCISION) & MULTS_6_1(52)(PERCISION downto 1))+signed(MULTS_6_2(52)(PERCISION) & MULTS_6_2(52)(PERCISION downto 1));
			MULTS_7_1(53)<=signed(MULTS_6_1(53)(PERCISION) & MULTS_6_1(53)(PERCISION downto 1))+signed(MULTS_6_2(53)(PERCISION) & MULTS_6_2(53)(PERCISION downto 1));
			MULTS_7_1(54)<=signed(MULTS_6_1(54)(PERCISION) & MULTS_6_1(54)(PERCISION downto 1))+signed(MULTS_6_2(54)(PERCISION) & MULTS_6_2(54)(PERCISION downto 1));
			MULTS_7_1(55)<=signed(MULTS_6_1(55)(PERCISION) & MULTS_6_1(55)(PERCISION downto 1))+signed(MULTS_6_2(55)(PERCISION) & MULTS_6_2(55)(PERCISION downto 1));
			MULTS_7_1(56)<=signed(MULTS_6_1(56)(PERCISION) & MULTS_6_1(56)(PERCISION downto 1))+signed(MULTS_6_2(56)(PERCISION) & MULTS_6_2(56)(PERCISION downto 1));
			MULTS_7_1(57)<=signed(MULTS_6_1(57)(PERCISION) & MULTS_6_1(57)(PERCISION downto 1))+signed(MULTS_6_2(57)(PERCISION) & MULTS_6_2(57)(PERCISION downto 1));
			MULTS_7_1(58)<=signed(MULTS_6_1(58)(PERCISION) & MULTS_6_1(58)(PERCISION downto 1))+signed(MULTS_6_2(58)(PERCISION) & MULTS_6_2(58)(PERCISION downto 1));
			MULTS_7_1(59)<=signed(MULTS_6_1(59)(PERCISION) & MULTS_6_1(59)(PERCISION downto 1))+signed(MULTS_6_2(59)(PERCISION) & MULTS_6_2(59)(PERCISION downto 1));
			MULTS_7_1(60)<=signed(MULTS_6_1(60)(PERCISION) & MULTS_6_1(60)(PERCISION downto 1))+signed(MULTS_6_2(60)(PERCISION) & MULTS_6_2(60)(PERCISION downto 1));
			MULTS_7_1(61)<=signed(MULTS_6_1(61)(PERCISION) & MULTS_6_1(61)(PERCISION downto 1))+signed(MULTS_6_2(61)(PERCISION) & MULTS_6_2(61)(PERCISION downto 1));
			MULTS_7_1(62)<=signed(MULTS_6_1(62)(PERCISION) & MULTS_6_1(62)(PERCISION downto 1))+signed(MULTS_6_2(62)(PERCISION) & MULTS_6_2(62)(PERCISION downto 1));
			MULTS_7_1(63)<=signed(MULTS_6_1(63)(PERCISION) & MULTS_6_1(63)(PERCISION downto 1))+signed(MULTS_6_2(63)(PERCISION) & MULTS_6_2(63)(PERCISION downto 1));
			MULTS_7_1(64)<=signed(MULTS_6_1(64)(PERCISION) & MULTS_6_1(64)(PERCISION downto 1))+signed(MULTS_6_2(64)(PERCISION) & MULTS_6_2(64)(PERCISION downto 1));
			MULTS_7_1(65)<=signed(MULTS_6_1(65)(PERCISION) & MULTS_6_1(65)(PERCISION downto 1))+signed(MULTS_6_2(65)(PERCISION) & MULTS_6_2(65)(PERCISION downto 1));
			MULTS_7_1(66)<=signed(MULTS_6_1(66)(PERCISION) & MULTS_6_1(66)(PERCISION downto 1))+signed(MULTS_6_2(66)(PERCISION) & MULTS_6_2(66)(PERCISION downto 1));
			MULTS_7_1(67)<=signed(MULTS_6_1(67)(PERCISION) & MULTS_6_1(67)(PERCISION downto 1))+signed(MULTS_6_2(67)(PERCISION) & MULTS_6_2(67)(PERCISION downto 1));
			MULTS_7_1(68)<=signed(MULTS_6_1(68)(PERCISION) & MULTS_6_1(68)(PERCISION downto 1))+signed(MULTS_6_2(68)(PERCISION) & MULTS_6_2(68)(PERCISION downto 1));
			MULTS_7_1(69)<=signed(MULTS_6_1(69)(PERCISION) & MULTS_6_1(69)(PERCISION downto 1))+signed(MULTS_6_2(69)(PERCISION) & MULTS_6_2(69)(PERCISION downto 1));
			MULTS_7_1(70)<=signed(MULTS_6_1(70)(PERCISION) & MULTS_6_1(70)(PERCISION downto 1))+signed(MULTS_6_2(70)(PERCISION) & MULTS_6_2(70)(PERCISION downto 1));
			MULTS_7_1(71)<=signed(MULTS_6_1(71)(PERCISION) & MULTS_6_1(71)(PERCISION downto 1))+signed(MULTS_6_2(71)(PERCISION) & MULTS_6_2(71)(PERCISION downto 1));
			MULTS_7_1(72)<=signed(MULTS_6_1(72)(PERCISION) & MULTS_6_1(72)(PERCISION downto 1))+signed(MULTS_6_2(72)(PERCISION) & MULTS_6_2(72)(PERCISION downto 1));
			MULTS_7_1(73)<=signed(MULTS_6_1(73)(PERCISION) & MULTS_6_1(73)(PERCISION downto 1))+signed(MULTS_6_2(73)(PERCISION) & MULTS_6_2(73)(PERCISION downto 1));
			MULTS_7_1(74)<=signed(MULTS_6_1(74)(PERCISION) & MULTS_6_1(74)(PERCISION downto 1))+signed(MULTS_6_2(74)(PERCISION) & MULTS_6_2(74)(PERCISION downto 1));
			MULTS_7_1(75)<=signed(MULTS_6_1(75)(PERCISION) & MULTS_6_1(75)(PERCISION downto 1))+signed(MULTS_6_2(75)(PERCISION) & MULTS_6_2(75)(PERCISION downto 1));
			MULTS_7_1(76)<=signed(MULTS_6_1(76)(PERCISION) & MULTS_6_1(76)(PERCISION downto 1))+signed(MULTS_6_2(76)(PERCISION) & MULTS_6_2(76)(PERCISION downto 1));
			MULTS_7_1(77)<=signed(MULTS_6_1(77)(PERCISION) & MULTS_6_1(77)(PERCISION downto 1))+signed(MULTS_6_2(77)(PERCISION) & MULTS_6_2(77)(PERCISION downto 1));
			MULTS_7_1(78)<=signed(MULTS_6_1(78)(PERCISION) & MULTS_6_1(78)(PERCISION downto 1))+signed(MULTS_6_2(78)(PERCISION) & MULTS_6_2(78)(PERCISION downto 1));
			MULTS_7_1(79)<=signed(MULTS_6_1(79)(PERCISION) & MULTS_6_1(79)(PERCISION downto 1))+signed(MULTS_6_2(79)(PERCISION) & MULTS_6_2(79)(PERCISION downto 1));
			MULTS_7_1(80)<=signed(MULTS_6_1(80)(PERCISION) & MULTS_6_1(80)(PERCISION downto 1))+signed(MULTS_6_2(80)(PERCISION) & MULTS_6_2(80)(PERCISION downto 1));
			MULTS_7_1(81)<=signed(MULTS_6_1(81)(PERCISION) & MULTS_6_1(81)(PERCISION downto 1))+signed(MULTS_6_2(81)(PERCISION) & MULTS_6_2(81)(PERCISION downto 1));
			MULTS_7_1(82)<=signed(MULTS_6_1(82)(PERCISION) & MULTS_6_1(82)(PERCISION downto 1))+signed(MULTS_6_2(82)(PERCISION) & MULTS_6_2(82)(PERCISION downto 1));
			MULTS_7_1(83)<=signed(MULTS_6_1(83)(PERCISION) & MULTS_6_1(83)(PERCISION downto 1))+signed(MULTS_6_2(83)(PERCISION) & MULTS_6_2(83)(PERCISION downto 1));



                        Enable_BIAS<='1';
		end if;


		------------------------------------STAGE-BIAS--------------------------------------
		if Enable_BIAS = '1' then

			BIAS_1<=(1+signed( MULTS_7_1(0)(PERCISION downto 1)));
			BIAS_2<=(1+signed( MULTS_7_1(1)(PERCISION downto 1)));
			BIAS_3<=(1+signed( MULTS_7_1(2)(PERCISION downto 1)));
			BIAS_4<=(1+signed( MULTS_7_1(3)(PERCISION downto 1)));
			BIAS_5<=(1+signed( MULTS_7_1(4)(PERCISION downto 1)));
			BIAS_6<=(1+signed( MULTS_7_1(5)(PERCISION downto 1)));
			BIAS_7<=(1+signed( MULTS_7_1(6)(PERCISION downto 1)));
			BIAS_8<=(1+signed( MULTS_7_1(7)(PERCISION downto 1)));
			BIAS_9<=(1+signed( MULTS_7_1(8)(PERCISION downto 1)));
			BIAS_10<=(1+signed( MULTS_7_1(9)(PERCISION downto 1)));
			BIAS_11<=(1+signed( MULTS_7_1(10)(PERCISION downto 1)));
			BIAS_12<=(1+signed( MULTS_7_1(11)(PERCISION downto 1)));
			BIAS_13<=(1+signed( MULTS_7_1(12)(PERCISION downto 1)));
			BIAS_14<=(1+signed( MULTS_7_1(13)(PERCISION downto 1)));
			BIAS_15<=(1+signed( MULTS_7_1(14)(PERCISION downto 1)));
			BIAS_16<=(1+signed( MULTS_7_1(15)(PERCISION downto 1)));
			BIAS_17<=(1+signed( MULTS_7_1(16)(PERCISION downto 1)));
			BIAS_18<=(1+signed( MULTS_7_1(17)(PERCISION downto 1)));
			BIAS_19<=(1+signed( MULTS_7_1(18)(PERCISION downto 1)));
			BIAS_20<=(1+signed( MULTS_7_1(19)(PERCISION downto 1)));
			BIAS_21<=(1+signed( MULTS_7_1(20)(PERCISION downto 1)));
			BIAS_22<=(1+signed( MULTS_7_1(21)(PERCISION downto 1)));
			BIAS_23<=(1+signed( MULTS_7_1(22)(PERCISION downto 1)));
			BIAS_24<=(1+signed( MULTS_7_1(23)(PERCISION downto 1)));
			BIAS_25<=(1+signed( MULTS_7_1(24)(PERCISION downto 1)));
			BIAS_26<=(1+signed( MULTS_7_1(25)(PERCISION downto 1)));
			BIAS_27<=(1+signed( MULTS_7_1(26)(PERCISION downto 1)));
			BIAS_28<=(1+signed( MULTS_7_1(27)(PERCISION downto 1)));
			BIAS_29<=(1+signed( MULTS_7_1(28)(PERCISION downto 1)));
			BIAS_30<=(1+signed( MULTS_7_1(29)(PERCISION downto 1)));
			BIAS_31<=(1+signed( MULTS_7_1(30)(PERCISION downto 1)));
			BIAS_32<=(1+signed( MULTS_7_1(31)(PERCISION downto 1)));
			BIAS_33<=(1+signed( MULTS_7_1(32)(PERCISION downto 1)));
			BIAS_34<=(1+signed( MULTS_7_1(33)(PERCISION downto 1)));
			BIAS_35<=(1+signed( MULTS_7_1(34)(PERCISION downto 1)));
			BIAS_36<=(1+signed( MULTS_7_1(35)(PERCISION downto 1)));
			BIAS_37<=(1+signed( MULTS_7_1(36)(PERCISION downto 1)));
			BIAS_38<=(1+signed( MULTS_7_1(37)(PERCISION downto 1)));
			BIAS_39<=(1+signed( MULTS_7_1(38)(PERCISION downto 1)));
			BIAS_40<=(1+signed( MULTS_7_1(39)(PERCISION downto 1)));
			BIAS_41<=(1+signed( MULTS_7_1(40)(PERCISION downto 1)));
			BIAS_42<=(1+signed( MULTS_7_1(41)(PERCISION downto 1)));
			BIAS_43<=(1+signed( MULTS_7_1(42)(PERCISION downto 1)));
			BIAS_44<=(1+signed( MULTS_7_1(43)(PERCISION downto 1)));
			BIAS_45<=(1+signed( MULTS_7_1(44)(PERCISION downto 1)));
			BIAS_46<=(1+signed( MULTS_7_1(45)(PERCISION downto 1)));
			BIAS_47<=(1+signed( MULTS_7_1(46)(PERCISION downto 1)));
			BIAS_48<=(1+signed( MULTS_7_1(47)(PERCISION downto 1)));
			BIAS_49<=(1+signed( MULTS_7_1(48)(PERCISION downto 1)));
			BIAS_50<=(1+signed( MULTS_7_1(49)(PERCISION downto 1)));
			BIAS_51<=(1+signed( MULTS_7_1(50)(PERCISION downto 1)));
			BIAS_52<=(1+signed( MULTS_7_1(51)(PERCISION downto 1)));
			BIAS_53<=(1+signed( MULTS_7_1(52)(PERCISION downto 1)));
			BIAS_54<=(1+signed( MULTS_7_1(53)(PERCISION downto 1)));
			BIAS_55<=(1+signed( MULTS_7_1(54)(PERCISION downto 1)));
			BIAS_56<=(1+signed( MULTS_7_1(55)(PERCISION downto 1)));
			BIAS_57<=(1+signed( MULTS_7_1(56)(PERCISION downto 1)));
			BIAS_58<=(1+signed( MULTS_7_1(57)(PERCISION downto 1)));
			BIAS_59<=(1+signed( MULTS_7_1(58)(PERCISION downto 1)));
			BIAS_60<=(1+signed( MULTS_7_1(59)(PERCISION downto 1)));
			BIAS_61<=(1+signed( MULTS_7_1(60)(PERCISION downto 1)));
			BIAS_62<=(1+signed( MULTS_7_1(61)(PERCISION downto 1)));
			BIAS_63<=(1+signed( MULTS_7_1(62)(PERCISION downto 1)));
			BIAS_64<=(1+signed( MULTS_7_1(63)(PERCISION downto 1)));
			BIAS_65<=(1+signed( MULTS_7_1(64)(PERCISION downto 1)));
			BIAS_66<=(1+signed( MULTS_7_1(65)(PERCISION downto 1)));
			BIAS_67<=(1+signed( MULTS_7_1(66)(PERCISION downto 1)));
			BIAS_68<=(1+signed( MULTS_7_1(67)(PERCISION downto 1)));
			BIAS_69<=(1+signed( MULTS_7_1(68)(PERCISION downto 1)));
			BIAS_70<=(1+signed( MULTS_7_1(69)(PERCISION downto 1)));
			BIAS_71<=(1+signed( MULTS_7_1(70)(PERCISION downto 1)));
			BIAS_72<=(1+signed( MULTS_7_1(71)(PERCISION downto 1)));
			BIAS_73<=(1+signed( MULTS_7_1(72)(PERCISION downto 1)));
			BIAS_74<=(1+signed( MULTS_7_1(73)(PERCISION downto 1)));
			BIAS_75<=(1+signed( MULTS_7_1(74)(PERCISION downto 1)));
			BIAS_76<=(1+signed( MULTS_7_1(75)(PERCISION downto 1)));
			BIAS_77<=(1+signed( MULTS_7_1(76)(PERCISION downto 1)));
			BIAS_78<=(1+signed( MULTS_7_1(77)(PERCISION downto 1)));
			BIAS_79<=(1+signed( MULTS_7_1(78)(PERCISION downto 1)));
			BIAS_80<=(1+signed( MULTS_7_1(79)(PERCISION downto 1)));
			BIAS_81<=(1+signed( MULTS_7_1(80)(PERCISION downto 1)));
			BIAS_82<=(1+signed( MULTS_7_1(81)(PERCISION downto 1)));
			BIAS_83<=(1+signed( MULTS_7_1(82)(PERCISION downto 1)));
			BIAS_84<=(1+signed( MULTS_7_1(83)(PERCISION downto 1)));

			Enable_ReLU<='1';
			
		end if;

		if SIG_STRIDE>1 and Enable_ReLU='1' then
                 SIG_STRIDE<=SIG_STRIDE-1; end if;

	if  Enable_ReLU='1' then
		if VALID_NXTLYR_PIX<VALID_LOCAL_PIX and SIG_STRIDE>(STRIDE-1) then

			if BIAS_1>0 then
			ReLU_1<=BIAS_1;
			DOUT_BUF_1_7<=std_logic_vector(BIAS_1);
			else
			ReLU_1<= (others => '0');
			DOUT_BUF_1_7<=(others => '0');
			end if;
			if BIAS_2>0 then
			ReLU_2<=BIAS_2;
			DOUT_BUF_2_7<=std_logic_vector(BIAS_2);
			else
			ReLU_2<= (others => '0');
			DOUT_BUF_2_7<=(others => '0');
			end if;
			if BIAS_3>0 then
			ReLU_3<=BIAS_3;
			DOUT_BUF_3_7<=std_logic_vector(BIAS_3);
			else
			ReLU_3<= (others => '0');
			DOUT_BUF_3_7<=(others => '0');
			end if;
			if BIAS_4>0 then
			ReLU_4<=BIAS_4;
			DOUT_BUF_4_7<=std_logic_vector(BIAS_4);
			else
			ReLU_4<= (others => '0');
			DOUT_BUF_4_7<=(others => '0');
			end if;
			if BIAS_5>0 then
			ReLU_5<=BIAS_5;
			DOUT_BUF_5_7<=std_logic_vector(BIAS_5);
			else
			ReLU_5<= (others => '0');
			DOUT_BUF_5_7<=(others => '0');
			end if;
			if BIAS_6>0 then
			ReLU_6<=BIAS_6;
			DOUT_BUF_6_7<=std_logic_vector(BIAS_6);
			else
			ReLU_6<= (others => '0');
			DOUT_BUF_6_7<=(others => '0');
			end if;
			if BIAS_7>0 then
			ReLU_7<=BIAS_7;
			DOUT_BUF_7_7<=std_logic_vector(BIAS_7);
			else
			ReLU_7<= (others => '0');
			DOUT_BUF_7_7<=(others => '0');
			end if;
			if BIAS_8>0 then
			ReLU_8<=BIAS_8;
			DOUT_BUF_8_7<=std_logic_vector(BIAS_8);
			else
			ReLU_8<= (others => '0');
			DOUT_BUF_8_7<=(others => '0');
			end if;
			if BIAS_9>0 then
			ReLU_9<=BIAS_9;
			DOUT_BUF_9_7<=std_logic_vector(BIAS_9);
			else
			ReLU_9<= (others => '0');
			DOUT_BUF_9_7<=(others => '0');
			end if;
			if BIAS_10>0 then
			ReLU_10<=BIAS_10;
			DOUT_BUF_10_7<=std_logic_vector(BIAS_10);
			else
			ReLU_10<= (others => '0');
			DOUT_BUF_10_7<=(others => '0');
			end if;
			if BIAS_11>0 then
			ReLU_11<=BIAS_11;
			DOUT_BUF_11_7<=std_logic_vector(BIAS_11);
			else
			ReLU_11<= (others => '0');
			DOUT_BUF_11_7<=(others => '0');
			end if;
			if BIAS_12>0 then
			ReLU_12<=BIAS_12;
			DOUT_BUF_12_7<=std_logic_vector(BIAS_12);
			else
			ReLU_12<= (others => '0');
			DOUT_BUF_12_7<=(others => '0');
			end if;
			if BIAS_13>0 then
			ReLU_13<=BIAS_13;
			DOUT_BUF_13_7<=std_logic_vector(BIAS_13);
			else
			ReLU_13<= (others => '0');
			DOUT_BUF_13_7<=(others => '0');
			end if;
			if BIAS_14>0 then
			ReLU_14<=BIAS_14;
			DOUT_BUF_14_7<=std_logic_vector(BIAS_14);
			else
			ReLU_14<= (others => '0');
			DOUT_BUF_14_7<=(others => '0');
			end if;
			if BIAS_15>0 then
			ReLU_15<=BIAS_15;
			DOUT_BUF_15_7<=std_logic_vector(BIAS_15);
			else
			ReLU_15<= (others => '0');
			DOUT_BUF_15_7<=(others => '0');
			end if;
			if BIAS_16>0 then
			ReLU_16<=BIAS_16;
			DOUT_BUF_16_7<=std_logic_vector(BIAS_16);
			else
			ReLU_16<= (others => '0');
			DOUT_BUF_16_7<=(others => '0');
			end if;
			if BIAS_17>0 then
			ReLU_17<=BIAS_17;
			DOUT_BUF_17_7<=std_logic_vector(BIAS_17);
			else
			ReLU_17<= (others => '0');
			DOUT_BUF_17_7<=(others => '0');
			end if;
			if BIAS_18>0 then
			ReLU_18<=BIAS_18;
			DOUT_BUF_18_7<=std_logic_vector(BIAS_18);
			else
			ReLU_18<= (others => '0');
			DOUT_BUF_18_7<=(others => '0');
			end if;
			if BIAS_19>0 then
			ReLU_19<=BIAS_19;
			DOUT_BUF_19_7<=std_logic_vector(BIAS_19);
			else
			ReLU_19<= (others => '0');
			DOUT_BUF_19_7<=(others => '0');
			end if;
			if BIAS_20>0 then
			ReLU_20<=BIAS_20;
			DOUT_BUF_20_7<=std_logic_vector(BIAS_20);
			else
			ReLU_20<= (others => '0');
			DOUT_BUF_20_7<=(others => '0');
			end if;
			if BIAS_21>0 then
			ReLU_21<=BIAS_21;
			DOUT_BUF_21_7<=std_logic_vector(BIAS_21);
			else
			ReLU_21<= (others => '0');
			DOUT_BUF_21_7<=(others => '0');
			end if;
			if BIAS_22>0 then
			ReLU_22<=BIAS_22;
			DOUT_BUF_22_7<=std_logic_vector(BIAS_22);
			else
			ReLU_22<= (others => '0');
			DOUT_BUF_22_7<=(others => '0');
			end if;
			if BIAS_23>0 then
			ReLU_23<=BIAS_23;
			DOUT_BUF_23_7<=std_logic_vector(BIAS_23);
			else
			ReLU_23<= (others => '0');
			DOUT_BUF_23_7<=(others => '0');
			end if;
			if BIAS_24>0 then
			ReLU_24<=BIAS_24;
			DOUT_BUF_24_7<=std_logic_vector(BIAS_24);
			else
			ReLU_24<= (others => '0');
			DOUT_BUF_24_7<=(others => '0');
			end if;
			if BIAS_25>0 then
			ReLU_25<=BIAS_25;
			DOUT_BUF_25_7<=std_logic_vector(BIAS_25);
			else
			ReLU_25<= (others => '0');
			DOUT_BUF_25_7<=(others => '0');
			end if;
			if BIAS_26>0 then
			ReLU_26<=BIAS_26;
			DOUT_BUF_26_7<=std_logic_vector(BIAS_26);
			else
			ReLU_26<= (others => '0');
			DOUT_BUF_26_7<=(others => '0');
			end if;
			if BIAS_27>0 then
			ReLU_27<=BIAS_27;
			DOUT_BUF_27_7<=std_logic_vector(BIAS_27);
			else
			ReLU_27<= (others => '0');
			DOUT_BUF_27_7<=(others => '0');
			end if;
			if BIAS_28>0 then
			ReLU_28<=BIAS_28;
			DOUT_BUF_28_7<=std_logic_vector(BIAS_28);
			else
			ReLU_28<= (others => '0');
			DOUT_BUF_28_7<=(others => '0');
			end if;
			if BIAS_29>0 then
			ReLU_29<=BIAS_29;
			DOUT_BUF_29_7<=std_logic_vector(BIAS_29);
			else
			ReLU_29<= (others => '0');
			DOUT_BUF_29_7<=(others => '0');
			end if;
			if BIAS_30>0 then
			ReLU_30<=BIAS_30;
			DOUT_BUF_30_7<=std_logic_vector(BIAS_30);
			else
			ReLU_30<= (others => '0');
			DOUT_BUF_30_7<=(others => '0');
			end if;
			if BIAS_31>0 then
			ReLU_31<=BIAS_31;
			DOUT_BUF_31_7<=std_logic_vector(BIAS_31);
			else
			ReLU_31<= (others => '0');
			DOUT_BUF_31_7<=(others => '0');
			end if;
			if BIAS_32>0 then
			ReLU_32<=BIAS_32;
			DOUT_BUF_32_7<=std_logic_vector(BIAS_32);
			else
			ReLU_32<= (others => '0');
			DOUT_BUF_32_7<=(others => '0');
			end if;
			if BIAS_33>0 then
			ReLU_33<=BIAS_33;
			DOUT_BUF_33_7<=std_logic_vector(BIAS_33);
			else
			ReLU_33<= (others => '0');
			DOUT_BUF_33_7<=(others => '0');
			end if;
			if BIAS_34>0 then
			ReLU_34<=BIAS_34;
			DOUT_BUF_34_7<=std_logic_vector(BIAS_34);
			else
			ReLU_34<= (others => '0');
			DOUT_BUF_34_7<=(others => '0');
			end if;
			if BIAS_35>0 then
			ReLU_35<=BIAS_35;
			DOUT_BUF_35_7<=std_logic_vector(BIAS_35);
			else
			ReLU_35<= (others => '0');
			DOUT_BUF_35_7<=(others => '0');
			end if;
			if BIAS_36>0 then
			ReLU_36<=BIAS_36;
			DOUT_BUF_36_7<=std_logic_vector(BIAS_36);
			else
			ReLU_36<= (others => '0');
			DOUT_BUF_36_7<=(others => '0');
			end if;
			if BIAS_37>0 then
			ReLU_37<=BIAS_37;
			DOUT_BUF_37_7<=std_logic_vector(BIAS_37);
			else
			ReLU_37<= (others => '0');
			DOUT_BUF_37_7<=(others => '0');
			end if;
			if BIAS_38>0 then
			ReLU_38<=BIAS_38;
			DOUT_BUF_38_7<=std_logic_vector(BIAS_38);
			else
			ReLU_38<= (others => '0');
			DOUT_BUF_38_7<=(others => '0');
			end if;
			if BIAS_39>0 then
			ReLU_39<=BIAS_39;
			DOUT_BUF_39_7<=std_logic_vector(BIAS_39);
			else
			ReLU_39<= (others => '0');
			DOUT_BUF_39_7<=(others => '0');
			end if;
			if BIAS_40>0 then
			ReLU_40<=BIAS_40;
			DOUT_BUF_40_7<=std_logic_vector(BIAS_40);
			else
			ReLU_40<= (others => '0');
			DOUT_BUF_40_7<=(others => '0');
			end if;
			if BIAS_41>0 then
			ReLU_41<=BIAS_41;
			DOUT_BUF_41_7<=std_logic_vector(BIAS_41);
			else
			ReLU_41<= (others => '0');
			DOUT_BUF_41_7<=(others => '0');
			end if;
			if BIAS_42>0 then
			ReLU_42<=BIAS_42;
			DOUT_BUF_42_7<=std_logic_vector(BIAS_42);
			else
			ReLU_42<= (others => '0');
			DOUT_BUF_42_7<=(others => '0');
			end if;
			if BIAS_43>0 then
			ReLU_43<=BIAS_43;
			DOUT_BUF_43_7<=std_logic_vector(BIAS_43);
			else
			ReLU_43<= (others => '0');
			DOUT_BUF_43_7<=(others => '0');
			end if;
			if BIAS_44>0 then
			ReLU_44<=BIAS_44;
			DOUT_BUF_44_7<=std_logic_vector(BIAS_44);
			else
			ReLU_44<= (others => '0');
			DOUT_BUF_44_7<=(others => '0');
			end if;
			if BIAS_45>0 then
			ReLU_45<=BIAS_45;
			DOUT_BUF_45_7<=std_logic_vector(BIAS_45);
			else
			ReLU_45<= (others => '0');
			DOUT_BUF_45_7<=(others => '0');
			end if;
			if BIAS_46>0 then
			ReLU_46<=BIAS_46;
			DOUT_BUF_46_7<=std_logic_vector(BIAS_46);
			else
			ReLU_46<= (others => '0');
			DOUT_BUF_46_7<=(others => '0');
			end if;
			if BIAS_47>0 then
			ReLU_47<=BIAS_47;
			DOUT_BUF_47_7<=std_logic_vector(BIAS_47);
			else
			ReLU_47<= (others => '0');
			DOUT_BUF_47_7<=(others => '0');
			end if;
			if BIAS_48>0 then
			ReLU_48<=BIAS_48;
			DOUT_BUF_48_7<=std_logic_vector(BIAS_48);
			else
			ReLU_48<= (others => '0');
			DOUT_BUF_48_7<=(others => '0');
			end if;
			if BIAS_49>0 then
			ReLU_49<=BIAS_49;
			DOUT_BUF_49_7<=std_logic_vector(BIAS_49);
			else
			ReLU_49<= (others => '0');
			DOUT_BUF_49_7<=(others => '0');
			end if;
			if BIAS_50>0 then
			ReLU_50<=BIAS_50;
			DOUT_BUF_50_7<=std_logic_vector(BIAS_50);
			else
			ReLU_50<= (others => '0');
			DOUT_BUF_50_7<=(others => '0');
			end if;
			if BIAS_51>0 then
			ReLU_51<=BIAS_51;
			DOUT_BUF_51_7<=std_logic_vector(BIAS_51);
			else
			ReLU_51<= (others => '0');
			DOUT_BUF_51_7<=(others => '0');
			end if;
			if BIAS_52>0 then
			ReLU_52<=BIAS_52;
			DOUT_BUF_52_7<=std_logic_vector(BIAS_52);
			else
			ReLU_52<= (others => '0');
			DOUT_BUF_52_7<=(others => '0');
			end if;
			if BIAS_53>0 then
			ReLU_53<=BIAS_53;
			DOUT_BUF_53_7<=std_logic_vector(BIAS_53);
			else
			ReLU_53<= (others => '0');
			DOUT_BUF_53_7<=(others => '0');
			end if;
			if BIAS_54>0 then
			ReLU_54<=BIAS_54;
			DOUT_BUF_54_7<=std_logic_vector(BIAS_54);
			else
			ReLU_54<= (others => '0');
			DOUT_BUF_54_7<=(others => '0');
			end if;
			if BIAS_55>0 then
			ReLU_55<=BIAS_55;
			DOUT_BUF_55_7<=std_logic_vector(BIAS_55);
			else
			ReLU_55<= (others => '0');
			DOUT_BUF_55_7<=(others => '0');
			end if;
			if BIAS_56>0 then
			ReLU_56<=BIAS_56;
			DOUT_BUF_56_7<=std_logic_vector(BIAS_56);
			else
			ReLU_56<= (others => '0');
			DOUT_BUF_56_7<=(others => '0');
			end if;
			if BIAS_57>0 then
			ReLU_57<=BIAS_57;
			DOUT_BUF_57_7<=std_logic_vector(BIAS_57);
			else
			ReLU_57<= (others => '0');
			DOUT_BUF_57_7<=(others => '0');
			end if;
			if BIAS_58>0 then
			ReLU_58<=BIAS_58;
			DOUT_BUF_58_7<=std_logic_vector(BIAS_58);
			else
			ReLU_58<= (others => '0');
			DOUT_BUF_58_7<=(others => '0');
			end if;
			if BIAS_59>0 then
			ReLU_59<=BIAS_59;
			DOUT_BUF_59_7<=std_logic_vector(BIAS_59);
			else
			ReLU_59<= (others => '0');
			DOUT_BUF_59_7<=(others => '0');
			end if;
			if BIAS_60>0 then
			ReLU_60<=BIAS_60;
			DOUT_BUF_60_7<=std_logic_vector(BIAS_60);
			else
			ReLU_60<= (others => '0');
			DOUT_BUF_60_7<=(others => '0');
			end if;
			if BIAS_61>0 then
			ReLU_61<=BIAS_61;
			DOUT_BUF_61_7<=std_logic_vector(BIAS_61);
			else
			ReLU_61<= (others => '0');
			DOUT_BUF_61_7<=(others => '0');
			end if;
			if BIAS_62>0 then
			ReLU_62<=BIAS_62;
			DOUT_BUF_62_7<=std_logic_vector(BIAS_62);
			else
			ReLU_62<= (others => '0');
			DOUT_BUF_62_7<=(others => '0');
			end if;
			if BIAS_63>0 then
			ReLU_63<=BIAS_63;
			DOUT_BUF_63_7<=std_logic_vector(BIAS_63);
			else
			ReLU_63<= (others => '0');
			DOUT_BUF_63_7<=(others => '0');
			end if;
			if BIAS_64>0 then
			ReLU_64<=BIAS_64;
			DOUT_BUF_64_7<=std_logic_vector(BIAS_64);
			else
			ReLU_64<= (others => '0');
			DOUT_BUF_64_7<=(others => '0');
			end if;
			if BIAS_65>0 then
			ReLU_65<=BIAS_65;
			DOUT_BUF_65_7<=std_logic_vector(BIAS_65);
			else
			ReLU_65<= (others => '0');
			DOUT_BUF_65_7<=(others => '0');
			end if;
			if BIAS_66>0 then
			ReLU_66<=BIAS_66;
			DOUT_BUF_66_7<=std_logic_vector(BIAS_66);
			else
			ReLU_66<= (others => '0');
			DOUT_BUF_66_7<=(others => '0');
			end if;
			if BIAS_67>0 then
			ReLU_67<=BIAS_67;
			DOUT_BUF_67_7<=std_logic_vector(BIAS_67);
			else
			ReLU_67<= (others => '0');
			DOUT_BUF_67_7<=(others => '0');
			end if;
			if BIAS_68>0 then
			ReLU_68<=BIAS_68;
			DOUT_BUF_68_7<=std_logic_vector(BIAS_68);
			else
			ReLU_68<= (others => '0');
			DOUT_BUF_68_7<=(others => '0');
			end if;
			if BIAS_69>0 then
			ReLU_69<=BIAS_69;
			DOUT_BUF_69_7<=std_logic_vector(BIAS_69);
			else
			ReLU_69<= (others => '0');
			DOUT_BUF_69_7<=(others => '0');
			end if;
			if BIAS_70>0 then
			ReLU_70<=BIAS_70;
			DOUT_BUF_70_7<=std_logic_vector(BIAS_70);
			else
			ReLU_70<= (others => '0');
			DOUT_BUF_70_7<=(others => '0');
			end if;
			if BIAS_71>0 then
			ReLU_71<=BIAS_71;
			DOUT_BUF_71_7<=std_logic_vector(BIAS_71);
			else
			ReLU_71<= (others => '0');
			DOUT_BUF_71_7<=(others => '0');
			end if;
			if BIAS_72>0 then
			ReLU_72<=BIAS_72;
			DOUT_BUF_72_7<=std_logic_vector(BIAS_72);
			else
			ReLU_72<= (others => '0');
			DOUT_BUF_72_7<=(others => '0');
			end if;
			if BIAS_73>0 then
			ReLU_73<=BIAS_73;
			DOUT_BUF_73_7<=std_logic_vector(BIAS_73);
			else
			ReLU_73<= (others => '0');
			DOUT_BUF_73_7<=(others => '0');
			end if;
			if BIAS_74>0 then
			ReLU_74<=BIAS_74;
			DOUT_BUF_74_7<=std_logic_vector(BIAS_74);
			else
			ReLU_74<= (others => '0');
			DOUT_BUF_74_7<=(others => '0');
			end if;
			if BIAS_75>0 then
			ReLU_75<=BIAS_75;
			DOUT_BUF_75_7<=std_logic_vector(BIAS_75);
			else
			ReLU_75<= (others => '0');
			DOUT_BUF_75_7<=(others => '0');
			end if;
			if BIAS_76>0 then
			ReLU_76<=BIAS_76;
			DOUT_BUF_76_7<=std_logic_vector(BIAS_76);
			else
			ReLU_76<= (others => '0');
			DOUT_BUF_76_7<=(others => '0');
			end if;
			if BIAS_77>0 then
			ReLU_77<=BIAS_77;
			DOUT_BUF_77_7<=std_logic_vector(BIAS_77);
			else
			ReLU_77<= (others => '0');
			DOUT_BUF_77_7<=(others => '0');
			end if;
			if BIAS_78>0 then
			ReLU_78<=BIAS_78;
			DOUT_BUF_78_7<=std_logic_vector(BIAS_78);
			else
			ReLU_78<= (others => '0');
			DOUT_BUF_78_7<=(others => '0');
			end if;
			if BIAS_79>0 then
			ReLU_79<=BIAS_79;
			DOUT_BUF_79_7<=std_logic_vector(BIAS_79);
			else
			ReLU_79<= (others => '0');
			DOUT_BUF_79_7<=(others => '0');
			end if;
			if BIAS_80>0 then
			ReLU_80<=BIAS_80;
			DOUT_BUF_80_7<=std_logic_vector(BIAS_80);
			else
			ReLU_80<= (others => '0');
			DOUT_BUF_80_7<=(others => '0');
			end if;
			if BIAS_81>0 then
			ReLU_81<=BIAS_81;
			DOUT_BUF_81_7<=std_logic_vector(BIAS_81);
			else
			ReLU_81<= (others => '0');
			DOUT_BUF_81_7<=(others => '0');
			end if;
			if BIAS_82>0 then
			ReLU_82<=BIAS_82;
			DOUT_BUF_82_7<=std_logic_vector(BIAS_82);
			else
			ReLU_82<= (others => '0');
			DOUT_BUF_82_7<=(others => '0');
			end if;
			if BIAS_83>0 then
			ReLU_83<=BIAS_83;
			DOUT_BUF_83_7<=std_logic_vector(BIAS_83);
			else
			ReLU_83<= (others => '0');
			DOUT_BUF_83_7<=(others => '0');
			end if;
			if BIAS_84>0 then
			ReLU_84<=BIAS_84;
			DOUT_BUF_84_7<=std_logic_vector(BIAS_84);
			else
			ReLU_84<= (others => '0');
			DOUT_BUF_84_7<=(others => '0');
			end if;

			EN_NXT_LYR_7<='1';FRST_TIM_EN_7<='1';
			OUT_PIXEL_COUNT<=OUT_PIXEL_COUNT+1;
		else
                       EN_NXT_LYR_7<='0';
                       DOUT_BUF_1_7<=(others => '0');
                       DOUT_BUF_2_7<=(others => '0');
                       DOUT_BUF_3_7<=(others => '0');
                       DOUT_BUF_4_7<=(others => '0');
                       DOUT_BUF_5_7<=(others => '0');
                       DOUT_BUF_6_7<=(others => '0');
                       DOUT_BUF_7_7<=(others => '0');
                       DOUT_BUF_8_7<=(others => '0');
                       DOUT_BUF_9_7<=(others => '0');
                       DOUT_BUF_10_7<=(others => '0');
                       DOUT_BUF_11_7<=(others => '0');
                       DOUT_BUF_12_7<=(others => '0');
                       DOUT_BUF_13_7<=(others => '0');
                       DOUT_BUF_14_7<=(others => '0');
                       DOUT_BUF_15_7<=(others => '0');
                       DOUT_BUF_16_7<=(others => '0');
                       DOUT_BUF_17_7<=(others => '0');
                       DOUT_BUF_18_7<=(others => '0');
                       DOUT_BUF_19_7<=(others => '0');
                       DOUT_BUF_20_7<=(others => '0');
                       DOUT_BUF_21_7<=(others => '0');
                       DOUT_BUF_22_7<=(others => '0');
                       DOUT_BUF_23_7<=(others => '0');
                       DOUT_BUF_24_7<=(others => '0');
                       DOUT_BUF_25_7<=(others => '0');
                       DOUT_BUF_26_7<=(others => '0');
                       DOUT_BUF_27_7<=(others => '0');
                       DOUT_BUF_28_7<=(others => '0');
                       DOUT_BUF_29_7<=(others => '0');
                       DOUT_BUF_30_7<=(others => '0');
                       DOUT_BUF_31_7<=(others => '0');
                       DOUT_BUF_32_7<=(others => '0');
                       DOUT_BUF_33_7<=(others => '0');
                       DOUT_BUF_34_7<=(others => '0');
                       DOUT_BUF_35_7<=(others => '0');
                       DOUT_BUF_36_7<=(others => '0');
                       DOUT_BUF_37_7<=(others => '0');
                       DOUT_BUF_38_7<=(others => '0');
                       DOUT_BUF_39_7<=(others => '0');
                       DOUT_BUF_40_7<=(others => '0');
                       DOUT_BUF_41_7<=(others => '0');
                       DOUT_BUF_42_7<=(others => '0');
                       DOUT_BUF_43_7<=(others => '0');
                       DOUT_BUF_44_7<=(others => '0');
                       DOUT_BUF_45_7<=(others => '0');
                       DOUT_BUF_46_7<=(others => '0');
                       DOUT_BUF_47_7<=(others => '0');
                       DOUT_BUF_48_7<=(others => '0');
                       DOUT_BUF_49_7<=(others => '0');
                       DOUT_BUF_50_7<=(others => '0');
                       DOUT_BUF_51_7<=(others => '0');
                       DOUT_BUF_52_7<=(others => '0');
                       DOUT_BUF_53_7<=(others => '0');
                       DOUT_BUF_54_7<=(others => '0');
                       DOUT_BUF_55_7<=(others => '0');
                       DOUT_BUF_56_7<=(others => '0');
                       DOUT_BUF_57_7<=(others => '0');
                       DOUT_BUF_58_7<=(others => '0');
                       DOUT_BUF_59_7<=(others => '0');
                       DOUT_BUF_60_7<=(others => '0');
                       DOUT_BUF_61_7<=(others => '0');
                       DOUT_BUF_62_7<=(others => '0');
                       DOUT_BUF_63_7<=(others => '0');
                       DOUT_BUF_64_7<=(others => '0');
                       DOUT_BUF_65_7<=(others => '0');
                       DOUT_BUF_66_7<=(others => '0');
                       DOUT_BUF_67_7<=(others => '0');
                       DOUT_BUF_68_7<=(others => '0');
                       DOUT_BUF_69_7<=(others => '0');
                       DOUT_BUF_70_7<=(others => '0');
                       DOUT_BUF_71_7<=(others => '0');
                       DOUT_BUF_72_7<=(others => '0');
                       DOUT_BUF_73_7<=(others => '0');
                       DOUT_BUF_74_7<=(others => '0');
                       DOUT_BUF_75_7<=(others => '0');
                       DOUT_BUF_76_7<=(others => '0');
                       DOUT_BUF_77_7<=(others => '0');
                       DOUT_BUF_78_7<=(others => '0');
                       DOUT_BUF_79_7<=(others => '0');
                       DOUT_BUF_80_7<=(others => '0');
                       DOUT_BUF_81_7<=(others => '0');
                       DOUT_BUF_82_7<=(others => '0');
                       DOUT_BUF_83_7<=(others => '0');
                       DOUT_BUF_84_7<=(others => '0');

		end if; -- VALIDPIXELS

		if VALID_NXTLYR_PIX=((VALID_LOCAL_PIX*STRIDE)-1) then VALID_NXTLYR_PIX<=0;SIG_STRIDE<=STRIDE;   -- reset sride and valid pixels
		else VALID_NXTLYR_PIX<=VALID_NXTLYR_PIX+1;end if; 

	end if;  --ReLU
elsif OUT_PIXEL_COUNT>=VALID_CYCLES  then INTERNAL_RST<='1';SIG_STRIDE<=STRIDE;EN_NXT_LYR_7<='1';  -- order is very important
else  EN_NXT_LYR_7<='0';-- In case stream stopped

end if; -- end enable 
end if; -- for RST	
end if; -- rising edge
end process LAYER_7;

EN_STREAM_OUT_7<= EN_STREAM_OUT_8;
VALID_OUT_7<= VALID_OUT_8;
DOUT_1_7<=DOUT_1_8;
DOUT_2_7<=DOUT_2_8;
DOUT_3_7<=DOUT_3_8;
DOUT_4_7<=DOUT_4_8;
DOUT_5_7<=DOUT_5_8;
DOUT_6_7<=DOUT_6_8;
DOUT_7_7<=DOUT_7_8;
DOUT_8_7<=DOUT_8_8;
DOUT_9_7<=DOUT_9_8;
DOUT_10_7<=DOUT_10_8;

end Behavioral;
------------------------------ ARCHITECTURE DECLARATION - END---------------------------------------------

