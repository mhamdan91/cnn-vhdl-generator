------------------------------------------HEADER START"------------------------------------------
--THIS FILE WAS GENERATED USING HIGH LANGUAGE DESCRIPTION TOOL DESIGNED BY: MUHAMMAD HAMDAN
--TOOL VERSION: 0.1
--GENERATION DATE/TIME:Mon Apr 06 09:41:57 CDT 2020
------------------------------------------HEADER END"--------------------------------------------



------------------------------DESCRIPTION AND LIBRARY DECLARATION-START---------------------------
-- Engineer:       Muhammad Hamdan
-- Design Name:    HDL GENERATION - CONV LAYER 
-- Module Name:    CONV - Behavioral 
-- Project Name:   CNN accelerator
-- Target Devices: Zynq-XC7Z020
-- Number of Total Operaiton: 832
-- Number of Clock Cycles: 11
-- Number of GOPS = 7.0
-- Description: 
-- Dependencies: 
-- Revision:0.010 


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_arith.all;

entity CONV_LAYER_3 is

GENERIC
 	( 
	constant PERCISION      : positive := 5; 	
	constant DOUT_WIDTH     : positive := 5; 	
	constant BIAS_SIZE      : positive := 5;	
	constant MULT_SIZE      : positive := 10;	
	constant DIN_WIDTH      : positive := 5;	
	constant IMAGE_WIDTH    : positive := 14;	
	constant IMAGE_SIZE     : positive := 1024;	
	constant F_SIZE         : positive := 5;	
	constant WEIGHT_SIZE    : positive := 5;	
	constant BIASES_SIZE	: positive := 2;
	constant PADDING        : positive := 1;	
	constant STRIDE         : positive := 1;	
	constant FEATURE_MAPS   : positive := 16;	
	constant VALID_CYCLES   : positive := 100;	
	constant STRIDE_CYCLES  : positive := 13;	
	constant VALID_LOCAL_PIX: positive := 10;	
	constant ADD_TREE_DEPTH : positive := 5;	
	constant INPUT_DEPTH    : positive := 3;
	constant FIFO_DEPTH     : positive := 10;	
	constant USED_FIFOS     : positive := 4;	
	constant MULT_SUM_D_1   : positive := 3;
	constant MULT_SUM_SIZE_1: positive := 6;
	constant MULT_SUM_D_2   : positive := 2;
	constant MULT_SUM_SIZE_2: positive := 6;
	constant MULT_SUM_D_3   : positive := 1;
	constant MULT_SUM_SIZE_3: positive := 6;
	constant ADD_1        : positive := 13;    	
	constant ADD_SIZE_1   : positive := 6;   	
	constant ADD_2        : positive := 7;    	
	constant ADD_SIZE_2   : positive := 6;   	
	constant ADD_3        : positive := 4;    	
	constant ADD_SIZE_3   : positive := 6;   	
	constant ADD_4        : positive := 2;    	
	constant ADD_SIZE_4   : positive := 6;   	
	constant ADD_5        : positive := 1;    	
	constant ADD_SIZE_5   : positive := 6;   	
	constant LOCAL_OUTPUT   : positive := 5	
		); 

port(
	DIN_1_3         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_2_3         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_3_3         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_4_3         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_5_3         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_6_3         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	CLK,RST         :IN std_logic;
   	DIS_STREAM      :OUT std_logic; 					-- S_AXIS_TVALID  : Data in is valid
   	EN_STREAM       :IN std_logic; 						-- S_AXIS_TREADY  : Ready to accept data in 
	EN_STREAM_OUT_3     :OUT std_logic; 				-- M_AXIS_TREADY  : Connected slave device is ready to accept data out/ Internal Enable
	VALID_OUT_3         :OUT std_logic;                             -- M_AXIS_TVALID  : Data out is valid
	EN_LOC_STREAM_3 :IN std_logic;
	DOUT_1_3            :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_2_3            :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_3_3            :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_4_3            :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_5_3            :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_6_3            :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_7_3            :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_8_3            :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_9_3            :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_10_3            :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	INTERNAL_RST        :OUT std_logic
	);	

end CONV_LAYER_3;

------------------------------ ARCHITECTURE DECLARATION - START---------------------------------------------

architecture Behavioral of CONV_LAYER_3 is

------------------------------ INTERNAL FIXED CONSTANT & SIGNALS DECLARATION - START---------------------------------------------
type       FILTER_TYPE             is array (0 to F_SIZE-1, 0 to F_SIZE-1) of signed(WEIGHT_SIZE- 1 downto 0);
type       FIFO_Memory             is array (0 to FIFO_DEPTH - 1)          of STD_LOGIC_VECTOR(DIN_WIDTH - 1 downto 0);
type       SLIDING_WINDOW          is array (0 to F_SIZE-1, 0 to F_SIZE-1) of STD_LOGIC_VECTOR(DIN_WIDTH- 1 downto 0);
signal     VALID_NXTLYR_PIX        :integer range 0 to STRIDE_CYCLES;
signal     PIXEL_COUNT             :integer range 0 to VALID_CYCLES;
signal     OUT_PIXEL_COUNT         :integer range 0 to VALID_CYCLES;
signal     EN_NXT_LYR_3            :std_logic;
signal     FRST_TIM_EN_3           :std_logic;
signal     Enable_MULT             :std_logic;
signal     Enable_ADDER            :std_logic;
signal     Enable_ReLU             :std_logic;
signal     Enable_BIAS             :std_logic;
signal     SIG_STRIDE              :integer range 0 to IMAGE_SIZE;
signal     PADDING_count           :integer range 0 to IMAGE_SIZE; -- TEMPORARY
signal     ROW_COUNT               :integer range 0 to IMAGE_SIZE; -- TEMPORARY
signal     WINDOW_1:SLIDING_WINDOW; 
signal     WINDOW_2:SLIDING_WINDOW; 
signal     WINDOW_3:SLIDING_WINDOW; 
signal     WINDOW_4:SLIDING_WINDOW; 
signal     WINDOW_5:SLIDING_WINDOW; 
signal     WINDOW_6:SLIDING_WINDOW; 


------------------------------ INTERNAL DYNAMIC SIGNALS DECLARATION ARRAY TYPE- START---------------------------------------------

type    AADD_DEPTH_1	is array (0 to ADD_1-1, 0 to FEATURE_MAPS-1 ) of signed(ADD_SIZE_1- 1 downto 0);
signal  ADD_DEPTH_1:AADD_DEPTH_1;
signal  Enable_STAGE_1	: std_logic;
type    AADD_DEPTH_2	is array (0 to ADD_2-1, 0 to FEATURE_MAPS-1 ) of signed(ADD_SIZE_2- 1 downto 0);
signal  ADD_DEPTH_2:AADD_DEPTH_2;
signal  Enable_STAGE_2	: std_logic;
type    AADD_DEPTH_3	is array (0 to ADD_3-1, 0 to FEATURE_MAPS-1 ) of signed(ADD_SIZE_3- 1 downto 0);
signal  ADD_DEPTH_3:AADD_DEPTH_3;
signal  Enable_STAGE_3	: std_logic;
type    AADD_DEPTH_4	is array (0 to ADD_4-1, 0 to FEATURE_MAPS-1 ) of signed(ADD_SIZE_4- 1 downto 0);
signal  ADD_DEPTH_4:AADD_DEPTH_4;
signal  Enable_STAGE_4	: std_logic;
type    AADD_DEPTH_5	is array (0 to ADD_5-1, 0 to FEATURE_MAPS-1 ) of signed(ADD_SIZE_5- 1 downto 0);
signal  ADD_DEPTH_5:AADD_DEPTH_5;
signal  Enable_STAGE_5	: std_logic;


------------------------------------------------------ MULT SUMMATION DECLARATION-----------------------------------------------------------
type    MULT_X_SUM_1	is array (0 to F_SIZE-1, 0 to F_SIZE-1 ) of signed(MULT_SUM_SIZE_1- 1 downto 0);
signal  EN_SUM_MULT_1	: std_logic;
signal  MULTS_1_1_1:MULT_X_SUM_1;
signal  MULTS_1_1_2:MULT_X_SUM_1;
signal  MULTS_1_1_3:MULT_X_SUM_1;
signal  MULTS_1_1_4:MULT_X_SUM_1;
signal  MULTS_1_1_5:MULT_X_SUM_1;
signal  MULTS_1_1_6:MULT_X_SUM_1;
signal  MULTS_1_2_1:MULT_X_SUM_1;
signal  MULTS_1_2_2:MULT_X_SUM_1;
signal  MULTS_1_2_3:MULT_X_SUM_1;
signal  MULTS_1_2_4:MULT_X_SUM_1;
signal  MULTS_1_2_5:MULT_X_SUM_1;
signal  MULTS_1_2_6:MULT_X_SUM_1;
signal  MULTS_1_3_1:MULT_X_SUM_1;
signal  MULTS_1_3_2:MULT_X_SUM_1;
signal  MULTS_1_3_3:MULT_X_SUM_1;
signal  MULTS_1_3_4:MULT_X_SUM_1;
signal  MULTS_1_3_5:MULT_X_SUM_1;
signal  MULTS_1_3_6:MULT_X_SUM_1;
signal  MULTS_1_4_1:MULT_X_SUM_1;
signal  MULTS_1_4_2:MULT_X_SUM_1;
signal  MULTS_1_4_3:MULT_X_SUM_1;
signal  MULTS_1_4_4:MULT_X_SUM_1;
signal  MULTS_1_4_5:MULT_X_SUM_1;
signal  MULTS_1_4_6:MULT_X_SUM_1;
signal  MULTS_1_5_1:MULT_X_SUM_1;
signal  MULTS_1_5_2:MULT_X_SUM_1;
signal  MULTS_1_5_3:MULT_X_SUM_1;
signal  MULTS_1_5_4:MULT_X_SUM_1;
signal  MULTS_1_5_5:MULT_X_SUM_1;
signal  MULTS_1_5_6:MULT_X_SUM_1;
signal  MULTS_1_6_1:MULT_X_SUM_1;
signal  MULTS_1_6_2:MULT_X_SUM_1;
signal  MULTS_1_6_3:MULT_X_SUM_1;
signal  MULTS_1_6_4:MULT_X_SUM_1;
signal  MULTS_1_6_5:MULT_X_SUM_1;
signal  MULTS_1_6_6:MULT_X_SUM_1;
signal  MULTS_1_7_1:MULT_X_SUM_1;
signal  MULTS_1_7_2:MULT_X_SUM_1;
signal  MULTS_1_7_3:MULT_X_SUM_1;
signal  MULTS_1_7_4:MULT_X_SUM_1;
signal  MULTS_1_7_5:MULT_X_SUM_1;
signal  MULTS_1_7_6:MULT_X_SUM_1;
signal  MULTS_1_8_1:MULT_X_SUM_1;
signal  MULTS_1_8_2:MULT_X_SUM_1;
signal  MULTS_1_8_3:MULT_X_SUM_1;
signal  MULTS_1_8_4:MULT_X_SUM_1;
signal  MULTS_1_8_5:MULT_X_SUM_1;
signal  MULTS_1_8_6:MULT_X_SUM_1;
signal  MULTS_1_9_1:MULT_X_SUM_1;
signal  MULTS_1_9_2:MULT_X_SUM_1;
signal  MULTS_1_9_3:MULT_X_SUM_1;
signal  MULTS_1_9_4:MULT_X_SUM_1;
signal  MULTS_1_9_5:MULT_X_SUM_1;
signal  MULTS_1_9_6:MULT_X_SUM_1;
signal  MULTS_1_10_1:MULT_X_SUM_1;
signal  MULTS_1_10_2:MULT_X_SUM_1;
signal  MULTS_1_10_3:MULT_X_SUM_1;
signal  MULTS_1_10_4:MULT_X_SUM_1;
signal  MULTS_1_10_5:MULT_X_SUM_1;
signal  MULTS_1_10_6:MULT_X_SUM_1;
signal  MULTS_1_11_1:MULT_X_SUM_1;
signal  MULTS_1_11_2:MULT_X_SUM_1;
signal  MULTS_1_11_3:MULT_X_SUM_1;
signal  MULTS_1_11_4:MULT_X_SUM_1;
signal  MULTS_1_11_5:MULT_X_SUM_1;
signal  MULTS_1_11_6:MULT_X_SUM_1;
signal  MULTS_1_12_1:MULT_X_SUM_1;
signal  MULTS_1_12_2:MULT_X_SUM_1;
signal  MULTS_1_12_3:MULT_X_SUM_1;
signal  MULTS_1_12_4:MULT_X_SUM_1;
signal  MULTS_1_12_5:MULT_X_SUM_1;
signal  MULTS_1_12_6:MULT_X_SUM_1;
signal  MULTS_1_13_1:MULT_X_SUM_1;
signal  MULTS_1_13_2:MULT_X_SUM_1;
signal  MULTS_1_13_3:MULT_X_SUM_1;
signal  MULTS_1_13_4:MULT_X_SUM_1;
signal  MULTS_1_13_5:MULT_X_SUM_1;
signal  MULTS_1_13_6:MULT_X_SUM_1;
signal  MULTS_1_14_1:MULT_X_SUM_1;
signal  MULTS_1_14_2:MULT_X_SUM_1;
signal  MULTS_1_14_3:MULT_X_SUM_1;
signal  MULTS_1_14_4:MULT_X_SUM_1;
signal  MULTS_1_14_5:MULT_X_SUM_1;
signal  MULTS_1_14_6:MULT_X_SUM_1;
signal  MULTS_1_15_1:MULT_X_SUM_1;
signal  MULTS_1_15_2:MULT_X_SUM_1;
signal  MULTS_1_15_3:MULT_X_SUM_1;
signal  MULTS_1_15_4:MULT_X_SUM_1;
signal  MULTS_1_15_5:MULT_X_SUM_1;
signal  MULTS_1_15_6:MULT_X_SUM_1;
signal  MULTS_1_16_1:MULT_X_SUM_1;
signal  MULTS_1_16_2:MULT_X_SUM_1;
signal  MULTS_1_16_3:MULT_X_SUM_1;
signal  MULTS_1_16_4:MULT_X_SUM_1;
signal  MULTS_1_16_5:MULT_X_SUM_1;
signal  MULTS_1_16_6:MULT_X_SUM_1;
type    MULT_X_SUM_2	is array (0 to F_SIZE-1, 0 to F_SIZE-1 ) of signed(MULT_SUM_SIZE_2- 1 downto 0);
signal  EN_SUM_MULT_2	: std_logic;
signal  MULTS_2_1_1:MULT_X_SUM_2;
signal  MULTS_2_1_2:MULT_X_SUM_2;
signal  MULTS_2_1_3:MULT_X_SUM_2;
signal  MULTS_2_1_4:MULT_X_SUM_2;
signal  MULTS_2_1_5:MULT_X_SUM_2;
signal  MULTS_2_1_6:MULT_X_SUM_2;
signal  MULTS_2_2_1:MULT_X_SUM_2;
signal  MULTS_2_2_2:MULT_X_SUM_2;
signal  MULTS_2_2_3:MULT_X_SUM_2;
signal  MULTS_2_2_4:MULT_X_SUM_2;
signal  MULTS_2_2_5:MULT_X_SUM_2;
signal  MULTS_2_2_6:MULT_X_SUM_2;
signal  MULTS_2_3_1:MULT_X_SUM_2;
signal  MULTS_2_3_2:MULT_X_SUM_2;
signal  MULTS_2_3_3:MULT_X_SUM_2;
signal  MULTS_2_3_4:MULT_X_SUM_2;
signal  MULTS_2_3_5:MULT_X_SUM_2;
signal  MULTS_2_3_6:MULT_X_SUM_2;
signal  MULTS_2_4_1:MULT_X_SUM_2;
signal  MULTS_2_4_2:MULT_X_SUM_2;
signal  MULTS_2_4_3:MULT_X_SUM_2;
signal  MULTS_2_4_4:MULT_X_SUM_2;
signal  MULTS_2_4_5:MULT_X_SUM_2;
signal  MULTS_2_4_6:MULT_X_SUM_2;
signal  MULTS_2_5_1:MULT_X_SUM_2;
signal  MULTS_2_5_2:MULT_X_SUM_2;
signal  MULTS_2_5_3:MULT_X_SUM_2;
signal  MULTS_2_5_4:MULT_X_SUM_2;
signal  MULTS_2_5_5:MULT_X_SUM_2;
signal  MULTS_2_5_6:MULT_X_SUM_2;
signal  MULTS_2_6_1:MULT_X_SUM_2;
signal  MULTS_2_6_2:MULT_X_SUM_2;
signal  MULTS_2_6_3:MULT_X_SUM_2;
signal  MULTS_2_6_4:MULT_X_SUM_2;
signal  MULTS_2_6_5:MULT_X_SUM_2;
signal  MULTS_2_6_6:MULT_X_SUM_2;
signal  MULTS_2_7_1:MULT_X_SUM_2;
signal  MULTS_2_7_2:MULT_X_SUM_2;
signal  MULTS_2_7_3:MULT_X_SUM_2;
signal  MULTS_2_7_4:MULT_X_SUM_2;
signal  MULTS_2_7_5:MULT_X_SUM_2;
signal  MULTS_2_7_6:MULT_X_SUM_2;
signal  MULTS_2_8_1:MULT_X_SUM_2;
signal  MULTS_2_8_2:MULT_X_SUM_2;
signal  MULTS_2_8_3:MULT_X_SUM_2;
signal  MULTS_2_8_4:MULT_X_SUM_2;
signal  MULTS_2_8_5:MULT_X_SUM_2;
signal  MULTS_2_8_6:MULT_X_SUM_2;
signal  MULTS_2_9_1:MULT_X_SUM_2;
signal  MULTS_2_9_2:MULT_X_SUM_2;
signal  MULTS_2_9_3:MULT_X_SUM_2;
signal  MULTS_2_9_4:MULT_X_SUM_2;
signal  MULTS_2_9_5:MULT_X_SUM_2;
signal  MULTS_2_9_6:MULT_X_SUM_2;
signal  MULTS_2_10_1:MULT_X_SUM_2;
signal  MULTS_2_10_2:MULT_X_SUM_2;
signal  MULTS_2_10_3:MULT_X_SUM_2;
signal  MULTS_2_10_4:MULT_X_SUM_2;
signal  MULTS_2_10_5:MULT_X_SUM_2;
signal  MULTS_2_10_6:MULT_X_SUM_2;
signal  MULTS_2_11_1:MULT_X_SUM_2;
signal  MULTS_2_11_2:MULT_X_SUM_2;
signal  MULTS_2_11_3:MULT_X_SUM_2;
signal  MULTS_2_11_4:MULT_X_SUM_2;
signal  MULTS_2_11_5:MULT_X_SUM_2;
signal  MULTS_2_11_6:MULT_X_SUM_2;
signal  MULTS_2_12_1:MULT_X_SUM_2;
signal  MULTS_2_12_2:MULT_X_SUM_2;
signal  MULTS_2_12_3:MULT_X_SUM_2;
signal  MULTS_2_12_4:MULT_X_SUM_2;
signal  MULTS_2_12_5:MULT_X_SUM_2;
signal  MULTS_2_12_6:MULT_X_SUM_2;
signal  MULTS_2_13_1:MULT_X_SUM_2;
signal  MULTS_2_13_2:MULT_X_SUM_2;
signal  MULTS_2_13_3:MULT_X_SUM_2;
signal  MULTS_2_13_4:MULT_X_SUM_2;
signal  MULTS_2_13_5:MULT_X_SUM_2;
signal  MULTS_2_13_6:MULT_X_SUM_2;
signal  MULTS_2_14_1:MULT_X_SUM_2;
signal  MULTS_2_14_2:MULT_X_SUM_2;
signal  MULTS_2_14_3:MULT_X_SUM_2;
signal  MULTS_2_14_4:MULT_X_SUM_2;
signal  MULTS_2_14_5:MULT_X_SUM_2;
signal  MULTS_2_14_6:MULT_X_SUM_2;
signal  MULTS_2_15_1:MULT_X_SUM_2;
signal  MULTS_2_15_2:MULT_X_SUM_2;
signal  MULTS_2_15_3:MULT_X_SUM_2;
signal  MULTS_2_15_4:MULT_X_SUM_2;
signal  MULTS_2_15_5:MULT_X_SUM_2;
signal  MULTS_2_15_6:MULT_X_SUM_2;
signal  MULTS_2_16_1:MULT_X_SUM_2;
signal  MULTS_2_16_2:MULT_X_SUM_2;
signal  MULTS_2_16_3:MULT_X_SUM_2;
signal  MULTS_2_16_4:MULT_X_SUM_2;
signal  MULTS_2_16_5:MULT_X_SUM_2;
signal  MULTS_2_16_6:MULT_X_SUM_2;
type    MULT_X_SUM_3	is array (0 to F_SIZE-1, 0 to F_SIZE-1 ) of signed(MULT_SUM_SIZE_3- 1 downto 0);
signal  EN_SUM_MULT_3	: std_logic;
signal  MULTS_3_1_1:MULT_X_SUM_3;
signal  MULTS_3_1_2:MULT_X_SUM_3;
signal  MULTS_3_1_3:MULT_X_SUM_3;
signal  MULTS_3_1_4:MULT_X_SUM_3;
signal  MULTS_3_1_5:MULT_X_SUM_3;
signal  MULTS_3_1_6:MULT_X_SUM_3;
signal  MULTS_3_2_1:MULT_X_SUM_3;
signal  MULTS_3_2_2:MULT_X_SUM_3;
signal  MULTS_3_2_3:MULT_X_SUM_3;
signal  MULTS_3_2_4:MULT_X_SUM_3;
signal  MULTS_3_2_5:MULT_X_SUM_3;
signal  MULTS_3_2_6:MULT_X_SUM_3;
signal  MULTS_3_3_1:MULT_X_SUM_3;
signal  MULTS_3_3_2:MULT_X_SUM_3;
signal  MULTS_3_3_3:MULT_X_SUM_3;
signal  MULTS_3_3_4:MULT_X_SUM_3;
signal  MULTS_3_3_5:MULT_X_SUM_3;
signal  MULTS_3_3_6:MULT_X_SUM_3;
signal  MULTS_3_4_1:MULT_X_SUM_3;
signal  MULTS_3_4_2:MULT_X_SUM_3;
signal  MULTS_3_4_3:MULT_X_SUM_3;
signal  MULTS_3_4_4:MULT_X_SUM_3;
signal  MULTS_3_4_5:MULT_X_SUM_3;
signal  MULTS_3_4_6:MULT_X_SUM_3;
signal  MULTS_3_5_1:MULT_X_SUM_3;
signal  MULTS_3_5_2:MULT_X_SUM_3;
signal  MULTS_3_5_3:MULT_X_SUM_3;
signal  MULTS_3_5_4:MULT_X_SUM_3;
signal  MULTS_3_5_5:MULT_X_SUM_3;
signal  MULTS_3_5_6:MULT_X_SUM_3;
signal  MULTS_3_6_1:MULT_X_SUM_3;
signal  MULTS_3_6_2:MULT_X_SUM_3;
signal  MULTS_3_6_3:MULT_X_SUM_3;
signal  MULTS_3_6_4:MULT_X_SUM_3;
signal  MULTS_3_6_5:MULT_X_SUM_3;
signal  MULTS_3_6_6:MULT_X_SUM_3;
signal  MULTS_3_7_1:MULT_X_SUM_3;
signal  MULTS_3_7_2:MULT_X_SUM_3;
signal  MULTS_3_7_3:MULT_X_SUM_3;
signal  MULTS_3_7_4:MULT_X_SUM_3;
signal  MULTS_3_7_5:MULT_X_SUM_3;
signal  MULTS_3_7_6:MULT_X_SUM_3;
signal  MULTS_3_8_1:MULT_X_SUM_3;
signal  MULTS_3_8_2:MULT_X_SUM_3;
signal  MULTS_3_8_3:MULT_X_SUM_3;
signal  MULTS_3_8_4:MULT_X_SUM_3;
signal  MULTS_3_8_5:MULT_X_SUM_3;
signal  MULTS_3_8_6:MULT_X_SUM_3;
signal  MULTS_3_9_1:MULT_X_SUM_3;
signal  MULTS_3_9_2:MULT_X_SUM_3;
signal  MULTS_3_9_3:MULT_X_SUM_3;
signal  MULTS_3_9_4:MULT_X_SUM_3;
signal  MULTS_3_9_5:MULT_X_SUM_3;
signal  MULTS_3_9_6:MULT_X_SUM_3;
signal  MULTS_3_10_1:MULT_X_SUM_3;
signal  MULTS_3_10_2:MULT_X_SUM_3;
signal  MULTS_3_10_3:MULT_X_SUM_3;
signal  MULTS_3_10_4:MULT_X_SUM_3;
signal  MULTS_3_10_5:MULT_X_SUM_3;
signal  MULTS_3_10_6:MULT_X_SUM_3;
signal  MULTS_3_11_1:MULT_X_SUM_3;
signal  MULTS_3_11_2:MULT_X_SUM_3;
signal  MULTS_3_11_3:MULT_X_SUM_3;
signal  MULTS_3_11_4:MULT_X_SUM_3;
signal  MULTS_3_11_5:MULT_X_SUM_3;
signal  MULTS_3_11_6:MULT_X_SUM_3;
signal  MULTS_3_12_1:MULT_X_SUM_3;
signal  MULTS_3_12_2:MULT_X_SUM_3;
signal  MULTS_3_12_3:MULT_X_SUM_3;
signal  MULTS_3_12_4:MULT_X_SUM_3;
signal  MULTS_3_12_5:MULT_X_SUM_3;
signal  MULTS_3_12_6:MULT_X_SUM_3;
signal  MULTS_3_13_1:MULT_X_SUM_3;
signal  MULTS_3_13_2:MULT_X_SUM_3;
signal  MULTS_3_13_3:MULT_X_SUM_3;
signal  MULTS_3_13_4:MULT_X_SUM_3;
signal  MULTS_3_13_5:MULT_X_SUM_3;
signal  MULTS_3_13_6:MULT_X_SUM_3;
signal  MULTS_3_14_1:MULT_X_SUM_3;
signal  MULTS_3_14_2:MULT_X_SUM_3;
signal  MULTS_3_14_3:MULT_X_SUM_3;
signal  MULTS_3_14_4:MULT_X_SUM_3;
signal  MULTS_3_14_5:MULT_X_SUM_3;
signal  MULTS_3_14_6:MULT_X_SUM_3;
signal  MULTS_3_15_1:MULT_X_SUM_3;
signal  MULTS_3_15_2:MULT_X_SUM_3;
signal  MULTS_3_15_3:MULT_X_SUM_3;
signal  MULTS_3_15_4:MULT_X_SUM_3;
signal  MULTS_3_15_5:MULT_X_SUM_3;
signal  MULTS_3_15_6:MULT_X_SUM_3;
signal  MULTS_3_16_1:MULT_X_SUM_3;
signal  MULTS_3_16_2:MULT_X_SUM_3;
signal  MULTS_3_16_3:MULT_X_SUM_3;
signal  MULTS_3_16_4:MULT_X_SUM_3;
signal  MULTS_3_16_5:MULT_X_SUM_3;
signal  MULTS_3_16_6:MULT_X_SUM_3;

type   MULT_X		is array (0 to F_SIZE-1, 0 to F_SIZE-1) of signed(MULT_SIZE-1 downto 0);
signal MULT_1_1:MULT_X;signal MULT_1_2:MULT_X;signal MULT_1_3:MULT_X;signal MULT_1_4:MULT_X;signal MULT_1_5:MULT_X;signal MULT_1_6:MULT_X;
signal DOUT_BUF_1_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_1		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_1		: signed(BIAS_SIZE-1   downto 0);

signal MULT_2_1:MULT_X;signal MULT_2_2:MULT_X;signal MULT_2_3:MULT_X;signal MULT_2_4:MULT_X;signal MULT_2_5:MULT_X;signal MULT_2_6:MULT_X;
signal DOUT_BUF_2_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_2		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_2		: signed(BIAS_SIZE-1   downto 0);

signal MULT_3_1:MULT_X;signal MULT_3_2:MULT_X;signal MULT_3_3:MULT_X;signal MULT_3_4:MULT_X;signal MULT_3_5:MULT_X;signal MULT_3_6:MULT_X;
signal DOUT_BUF_3_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_3		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_3		: signed(BIAS_SIZE-1   downto 0);

signal MULT_4_1:MULT_X;signal MULT_4_2:MULT_X;signal MULT_4_3:MULT_X;signal MULT_4_4:MULT_X;signal MULT_4_5:MULT_X;signal MULT_4_6:MULT_X;
signal DOUT_BUF_4_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_4		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_4		: signed(BIAS_SIZE-1   downto 0);

signal MULT_5_1:MULT_X;signal MULT_5_2:MULT_X;signal MULT_5_3:MULT_X;signal MULT_5_4:MULT_X;signal MULT_5_5:MULT_X;signal MULT_5_6:MULT_X;
signal DOUT_BUF_5_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_5		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_5		: signed(BIAS_SIZE-1   downto 0);

signal MULT_6_1:MULT_X;signal MULT_6_2:MULT_X;signal MULT_6_3:MULT_X;signal MULT_6_4:MULT_X;signal MULT_6_5:MULT_X;signal MULT_6_6:MULT_X;
signal DOUT_BUF_6_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_6		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_6		: signed(BIAS_SIZE-1   downto 0);

signal MULT_7_1:MULT_X;signal MULT_7_2:MULT_X;signal MULT_7_3:MULT_X;signal MULT_7_4:MULT_X;signal MULT_7_5:MULT_X;signal MULT_7_6:MULT_X;
signal DOUT_BUF_7_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_7		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_7		: signed(BIAS_SIZE-1   downto 0);

signal MULT_8_1:MULT_X;signal MULT_8_2:MULT_X;signal MULT_8_3:MULT_X;signal MULT_8_4:MULT_X;signal MULT_8_5:MULT_X;signal MULT_8_6:MULT_X;
signal DOUT_BUF_8_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_8		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_8		: signed(BIAS_SIZE-1   downto 0);

signal MULT_9_1:MULT_X;signal MULT_9_2:MULT_X;signal MULT_9_3:MULT_X;signal MULT_9_4:MULT_X;signal MULT_9_5:MULT_X;signal MULT_9_6:MULT_X;
signal DOUT_BUF_9_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_9		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_9		: signed(BIAS_SIZE-1   downto 0);

signal MULT_10_1:MULT_X;signal MULT_10_2:MULT_X;signal MULT_10_3:MULT_X;signal MULT_10_4:MULT_X;signal MULT_10_5:MULT_X;signal MULT_10_6:MULT_X;
signal DOUT_BUF_10_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_10		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_10		: signed(BIAS_SIZE-1   downto 0);

signal MULT_11_1:MULT_X;signal MULT_11_2:MULT_X;signal MULT_11_3:MULT_X;signal MULT_11_4:MULT_X;signal MULT_11_5:MULT_X;signal MULT_11_6:MULT_X;
signal DOUT_BUF_11_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_11		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_11		: signed(BIAS_SIZE-1   downto 0);

signal MULT_12_1:MULT_X;signal MULT_12_2:MULT_X;signal MULT_12_3:MULT_X;signal MULT_12_4:MULT_X;signal MULT_12_5:MULT_X;signal MULT_12_6:MULT_X;
signal DOUT_BUF_12_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_12		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_12		: signed(BIAS_SIZE-1   downto 0);

signal MULT_13_1:MULT_X;signal MULT_13_2:MULT_X;signal MULT_13_3:MULT_X;signal MULT_13_4:MULT_X;signal MULT_13_5:MULT_X;signal MULT_13_6:MULT_X;
signal DOUT_BUF_13_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_13		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_13		: signed(BIAS_SIZE-1   downto 0);

signal MULT_14_1:MULT_X;signal MULT_14_2:MULT_X;signal MULT_14_3:MULT_X;signal MULT_14_4:MULT_X;signal MULT_14_5:MULT_X;signal MULT_14_6:MULT_X;
signal DOUT_BUF_14_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_14		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_14		: signed(BIAS_SIZE-1   downto 0);

signal MULT_15_1:MULT_X;signal MULT_15_2:MULT_X;signal MULT_15_3:MULT_X;signal MULT_15_4:MULT_X;signal MULT_15_5:MULT_X;signal MULT_15_6:MULT_X;
signal DOUT_BUF_15_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_15		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_15		: signed(BIAS_SIZE-1   downto 0);

signal MULT_16_1:MULT_X;signal MULT_16_2:MULT_X;signal MULT_16_3:MULT_X;signal MULT_16_4:MULT_X;signal MULT_16_5:MULT_X;signal MULT_16_6:MULT_X;
signal DOUT_BUF_16_3	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_16		: signed(BIAS_SIZE-1   downto 0);
signal ReLU_16		: signed(BIAS_SIZE-1   downto 0);



------------------------------------------------------ FIFO_1_1 DECLARATION---------------------------------------------------------
signal FIFO_1_ROW_1  	: FIFO_Memory;
signal HEAD_1_1       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_1_1       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_1_1	: std_logic;
signal ReadEn_1_1 	: std_logic;
signal Async_Mode_1_1 : boolean;

------------------------------------------------------ FIFO_2_1 DECLARATION---------------------------------------------------------
signal FIFO_2_ROW_1  	: FIFO_Memory;
signal HEAD_2_1       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_2_1       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_2_1	: std_logic;
signal ReadEn_2_1 	: std_logic;
signal Async_Mode_2_1 : boolean;

------------------------------------------------------ FIFO_3_1 DECLARATION---------------------------------------------------------
signal FIFO_3_ROW_1  	: FIFO_Memory;
signal HEAD_3_1       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_3_1       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_3_1	: std_logic;
signal ReadEn_3_1 	: std_logic;
signal Async_Mode_3_1 : boolean;

------------------------------------------------------ FIFO_4_1 DECLARATION---------------------------------------------------------
signal FIFO_4_ROW_1  	: FIFO_Memory;
signal HEAD_4_1       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_4_1       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_4_1	: std_logic;
signal ReadEn_4_1 	: std_logic;
signal Async_Mode_4_1 : boolean;

------------------------------------------------------ FIFO_5_1 DECLARATION---------------------------------------------------------
signal FIFO_5_ROW_1  	: FIFO_Memory;
signal HEAD_5_1       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_5_1       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_5_1	: std_logic;
signal ReadEn_5_1 	: std_logic;
signal Async_Mode_5_1 : boolean;

------------------------------------------------------ FIFO_6_1 DECLARATION---------------------------------------------------------
signal FIFO_6_ROW_1  	: FIFO_Memory;
signal HEAD_6_1       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_6_1       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_6_1	: std_logic;
signal ReadEn_6_1 	: std_logic;
signal Async_Mode_6_1 : boolean;

------------------------------------------------------ FIFO_1_2 DECLARATION---------------------------------------------------------
signal FIFO_1_ROW_2  	: FIFO_Memory;
signal HEAD_1_2       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_1_2       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_1_2	: std_logic;
signal ReadEn_1_2 	: std_logic;
signal Async_Mode_1_2 : boolean;

------------------------------------------------------ FIFO_2_2 DECLARATION---------------------------------------------------------
signal FIFO_2_ROW_2  	: FIFO_Memory;
signal HEAD_2_2       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_2_2       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_2_2	: std_logic;
signal ReadEn_2_2 	: std_logic;
signal Async_Mode_2_2 : boolean;

------------------------------------------------------ FIFO_3_2 DECLARATION---------------------------------------------------------
signal FIFO_3_ROW_2  	: FIFO_Memory;
signal HEAD_3_2       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_3_2       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_3_2	: std_logic;
signal ReadEn_3_2 	: std_logic;
signal Async_Mode_3_2 : boolean;

------------------------------------------------------ FIFO_4_2 DECLARATION---------------------------------------------------------
signal FIFO_4_ROW_2  	: FIFO_Memory;
signal HEAD_4_2       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_4_2       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_4_2	: std_logic;
signal ReadEn_4_2 	: std_logic;
signal Async_Mode_4_2 : boolean;

------------------------------------------------------ FIFO_5_2 DECLARATION---------------------------------------------------------
signal FIFO_5_ROW_2  	: FIFO_Memory;
signal HEAD_5_2       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_5_2       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_5_2	: std_logic;
signal ReadEn_5_2 	: std_logic;
signal Async_Mode_5_2 : boolean;

------------------------------------------------------ FIFO_6_2 DECLARATION---------------------------------------------------------
signal FIFO_6_ROW_2  	: FIFO_Memory;
signal HEAD_6_2       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_6_2       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_6_2	: std_logic;
signal ReadEn_6_2 	: std_logic;
signal Async_Mode_6_2 : boolean;

------------------------------------------------------ FIFO_1_3 DECLARATION---------------------------------------------------------
signal FIFO_1_ROW_3  	: FIFO_Memory;
signal HEAD_1_3       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_1_3       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_1_3	: std_logic;
signal ReadEn_1_3 	: std_logic;
signal Async_Mode_1_3 : boolean;

------------------------------------------------------ FIFO_2_3 DECLARATION---------------------------------------------------------
signal FIFO_2_ROW_3  	: FIFO_Memory;
signal HEAD_2_3       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_2_3       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_2_3	: std_logic;
signal ReadEn_2_3 	: std_logic;
signal Async_Mode_2_3 : boolean;

------------------------------------------------------ FIFO_3_3 DECLARATION---------------------------------------------------------
signal FIFO_3_ROW_3  	: FIFO_Memory;
signal HEAD_3_3       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_3_3       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_3_3	: std_logic;
signal ReadEn_3_3 	: std_logic;
signal Async_Mode_3_3 : boolean;

------------------------------------------------------ FIFO_4_3 DECLARATION---------------------------------------------------------
signal FIFO_4_ROW_3  	: FIFO_Memory;
signal HEAD_4_3       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_4_3       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_4_3	: std_logic;
signal ReadEn_4_3 	: std_logic;
signal Async_Mode_4_3 : boolean;

------------------------------------------------------ FIFO_5_3 DECLARATION---------------------------------------------------------
signal FIFO_5_ROW_3  	: FIFO_Memory;
signal HEAD_5_3       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_5_3       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_5_3	: std_logic;
signal ReadEn_5_3 	: std_logic;
signal Async_Mode_5_3 : boolean;

------------------------------------------------------ FIFO_6_3 DECLARATION---------------------------------------------------------
signal FIFO_6_ROW_3  	: FIFO_Memory;
signal HEAD_6_3       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_6_3       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_6_3	: std_logic;
signal ReadEn_6_3 	: std_logic;
signal Async_Mode_6_3 : boolean;

------------------------------------------------------ FIFO_1_4 DECLARATION---------------------------------------------------------
signal FIFO_1_ROW_4  	: FIFO_Memory;
signal HEAD_1_4       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_1_4       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_1_4	: std_logic;
signal ReadEn_1_4 	: std_logic;
signal Async_Mode_1_4 : boolean;

------------------------------------------------------ FIFO_2_4 DECLARATION---------------------------------------------------------
signal FIFO_2_ROW_4  	: FIFO_Memory;
signal HEAD_2_4       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_2_4       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_2_4	: std_logic;
signal ReadEn_2_4 	: std_logic;
signal Async_Mode_2_4 : boolean;

------------------------------------------------------ FIFO_3_4 DECLARATION---------------------------------------------------------
signal FIFO_3_ROW_4  	: FIFO_Memory;
signal HEAD_3_4       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_3_4       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_3_4	: std_logic;
signal ReadEn_3_4 	: std_logic;
signal Async_Mode_3_4 : boolean;

------------------------------------------------------ FIFO_4_4 DECLARATION---------------------------------------------------------
signal FIFO_4_ROW_4  	: FIFO_Memory;
signal HEAD_4_4       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_4_4       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_4_4	: std_logic;
signal ReadEn_4_4 	: std_logic;
signal Async_Mode_4_4 : boolean;

------------------------------------------------------ FIFO_5_4 DECLARATION---------------------------------------------------------
signal FIFO_5_ROW_4  	: FIFO_Memory;
signal HEAD_5_4       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_5_4       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_5_4	: std_logic;
signal ReadEn_5_4 	: std_logic;
signal Async_Mode_5_4 : boolean;

------------------------------------------------------ FIFO_6_4 DECLARATION---------------------------------------------------------
signal FIFO_6_ROW_4  	: FIFO_Memory;
signal HEAD_6_4       : natural range 0 to FIFO_DEPTH - 1;
signal TAIL_6_4       : natural range 0 to FIFO_DEPTH - 1;
signal WriteEn_6_4	: std_logic;
signal ReadEn_6_4 	: std_logic;
signal Async_Mode_6_4 : boolean;


-------------------------------------- OUTPUT FROM LOWER COMPONENT SIGNALS--------------------------------------------------
signal DOUT_1_4          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_2_4          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_3_4          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_4_4          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_5_4          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_6_4          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_7_4          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_8_4          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_9_4          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal DOUT_10_4          : std_logic_vector(DOUT_WIDTH-1 downto 0);
signal EN_STREAM_OUT_4	 : std_logic;
signal VALID_OUT_4       : std_logic;

--------------------------------------------- FILTER HARDCODED CONSTANTS -WEIGHTS START--------------------------------

constant FMAP_1_1: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_1: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_1: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_1: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_1: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_1: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_2: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_2: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_2: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_2: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_2: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_2: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_3: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_3: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_3: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_3: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_3: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_3: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_4: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_4: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_4: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_4: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_4: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_4: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_5: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_5: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_5: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_5: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_5: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_5: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_6: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_6: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_6: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_6: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_6: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_6: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_7: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_7: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_7: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_7: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_7: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_7: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_8: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_8: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_8: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_8: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_8: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_8: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_9: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_9: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_9: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_9: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_9: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_9: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_10: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_10: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_10: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_10: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_10: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_10: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_11: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_11: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_11: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_11: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_11: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_11: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_12: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_12: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_12: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_12: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_12: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_12: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_13: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_13: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_13: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_13: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_13: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_13: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_14: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_14: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_14: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_14: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_14: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_14: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_15: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_15: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_15: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_15: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_15: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_15: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_1_16: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_2_16: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_3_16: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_4_16: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_5_16: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );

constant FMAP_6_16: FILTER_TYPE:=		(("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001"),
                                     ("00001","00010","00011","00010","00001")
                                    );


constant BIAS_VAL_1: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_2: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_3: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_4: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_5: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_6: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_7: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_8: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_9: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_10: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_11: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_12: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_13: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_14: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_15: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_16: signed (BIASES_SIZE-1 downto 0):="01";


---------------------------------- MAP NEXT LAYER - COMPONENTS START----------------------------------
COMPONENT POOL_LAYER_4
    port(	CLK,RST			:IN std_logic;
		DIN_1_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_2_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_3_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_4_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_5_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_6_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_7_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_8_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_9_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_10_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_11_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_12_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_13_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_14_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_15_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		DIN_16_4		:IN std_logic_vector(LOCAL_OUTPUT-1 downto 0);
		EN_STREAM_OUT_4	:OUT std_logic;
		VALID_OUT_4		:OUT std_logic;
		DOUT_1_4        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_2_4        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_3_4        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_4_4        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_5_4        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_6_4        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_7_4        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_8_4        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_9_4        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		DOUT_10_4        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
		EN_STREAM		:IN std_logic;
		EN_LOC_STREAM_4	:IN std_logic
      			);
END COMPONENT POOL_LAYER_4;

begin

POOL_LYR_4 : POOL_LAYER_4 
          port map(
          CLK                 => CLK,
          RST                 => RST,
          DIN_1_4             => DOUT_BUF_1_3,
          DIN_2_4             => DOUT_BUF_2_3,
          DIN_3_4             => DOUT_BUF_3_3,
          DIN_4_4             => DOUT_BUF_4_3,
          DIN_5_4             => DOUT_BUF_5_3,
          DIN_6_4             => DOUT_BUF_6_3,
          DIN_7_4             => DOUT_BUF_7_3,
          DIN_8_4             => DOUT_BUF_8_3,
          DIN_9_4             => DOUT_BUF_9_3,
          DIN_10_4             => DOUT_BUF_10_3,
          DIN_11_4             => DOUT_BUF_11_3,
          DIN_12_4             => DOUT_BUF_12_3,
          DIN_13_4             => DOUT_BUF_13_3,
          DIN_14_4             => DOUT_BUF_14_3,
          DIN_15_4             => DOUT_BUF_15_3,
          DIN_16_4             => DOUT_BUF_16_3,
          DOUT_1_4            => DOUT_1_4,
          DOUT_2_4            => DOUT_2_4,
          DOUT_3_4            => DOUT_3_4,
          DOUT_4_4            => DOUT_4_4,
          DOUT_5_4            => DOUT_5_4,
          DOUT_6_4            => DOUT_6_4,
          DOUT_7_4            => DOUT_7_4,
          DOUT_8_4            => DOUT_8_4,
          DOUT_9_4            => DOUT_9_4,
          DOUT_10_4            => DOUT_10_4,
          VALID_OUT_4         => VALID_OUT_4,
          EN_STREAM_OUT_4     => EN_STREAM_OUT_4,
          EN_LOC_STREAM_4     => EN_NXT_LYR_3,
          EN_STREAM           => EN_STREAM
                );

----------------------------------------------- MAP NEXT LAYER - COMPONENTS END----------------------------------------------------



-------------------------------------------------------- ARCHITECTURE BEGIN--------------------------------------------------------

LAYER_3: process(CLK)


begin
------------------------------------------------ RESET AND PROCESS TOP START ------------------------------------------------------
if rising_edge(CLK) then
  if RST = '1' then
	-------------------FIXED SIGNALS RESET------------------------
    PIXEL_COUNT<=0;VALID_NXTLYR_PIX<=0;OUT_PIXEL_COUNT<=0;
    EN_NXT_LYR_3<='0';FRST_TIM_EN_3<='0';
    Enable_MULT<='0';Enable_ADDER<='0';Enable_ReLU<='0';Enable_BIAS<='0';
    INTERNAL_RST<='0';PADDING_count<=0;ROW_COUNT<=0;SIG_STRIDE<=STRIDE;

-------------------DYNAMIC SIGNALS RESET------------------------
    WINDOW_1<=((others=> (others=> (others=>'0'))));
    WINDOW_2<=((others=> (others=> (others=>'0'))));
    WINDOW_3<=((others=> (others=> (others=>'0'))));
    WINDOW_4<=((others=> (others=> (others=>'0'))));
    WINDOW_5<=((others=> (others=> (others=>'0'))));
    WINDOW_6<=((others=> (others=> (others=>'0'))));

    MULTS_1_1_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_6<=((others=> (others=> (others=>'0'))));
    EN_SUM_MULT_1<='0';
    MULTS_1_1_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_1_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_1_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_1_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_1_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_1_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_1_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_2_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_2_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_2_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_2_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_2_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_2_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_3_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_3_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_3_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_3_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_3_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_3_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_4_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_4_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_4_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_4_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_4_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_4_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_5_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_5_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_5_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_5_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_5_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_5_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_6_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_6_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_6_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_6_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_6_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_6_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_7_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_7_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_7_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_7_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_7_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_7_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_8_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_8_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_8_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_8_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_8_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_8_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_9_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_9_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_9_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_9_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_9_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_9_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_10_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_10_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_10_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_10_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_10_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_10_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_11_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_11_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_11_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_11_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_11_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_11_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_12_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_12_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_12_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_12_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_12_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_12_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_13_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_13_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_13_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_13_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_13_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_13_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_14_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_14_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_14_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_14_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_14_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_14_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_15_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_15_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_15_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_15_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_15_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_15_6<=((others=> (others=> (others=>'0'))));
    EN_SUM_MULT_2<='0';
    MULTS_1_1_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_1_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_2_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_3_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_4_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_5_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_6_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_7_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_8_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_9_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_10_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_11_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_12_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_13_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_14_6<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_1<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_2<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_3<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_4<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_5<=((others=> (others=> (others=>'0'))));
    MULTS_1_15_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_1_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_1_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_1_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_1_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_1_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_1_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_2_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_2_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_2_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_2_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_2_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_2_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_3_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_3_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_3_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_3_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_3_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_3_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_4_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_4_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_4_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_4_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_4_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_4_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_5_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_5_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_5_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_5_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_5_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_5_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_6_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_6_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_6_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_6_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_6_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_6_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_7_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_7_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_7_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_7_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_7_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_7_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_8_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_8_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_8_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_8_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_8_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_8_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_9_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_9_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_9_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_9_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_9_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_9_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_10_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_10_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_10_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_10_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_10_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_10_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_11_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_11_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_11_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_11_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_11_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_11_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_12_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_12_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_12_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_12_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_12_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_12_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_13_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_13_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_13_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_13_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_13_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_13_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_14_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_14_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_14_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_14_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_14_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_14_6<=((others=> (others=> (others=>'0'))));
    MULTS_2_15_1<=((others=> (others=> (others=>'0'))));
    MULTS_2_15_2<=((others=> (others=> (others=>'0'))));
    MULTS_2_15_3<=((others=> (others=> (others=>'0'))));
    MULTS_2_15_4<=((others=> (others=> (others=>'0'))));
    MULTS_2_15_5<=((others=> (others=> (others=>'0'))));
    MULTS_2_15_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_1_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_1_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_1_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_1_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_1_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_1_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_2_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_2_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_2_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_2_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_2_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_2_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_3_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_3_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_3_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_3_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_3_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_3_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_4_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_4_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_4_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_4_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_4_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_4_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_5_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_5_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_5_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_5_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_5_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_5_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_6_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_6_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_6_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_6_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_6_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_6_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_7_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_7_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_7_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_7_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_7_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_7_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_8_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_8_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_8_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_8_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_8_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_8_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_9_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_9_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_9_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_9_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_9_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_9_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_10_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_10_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_10_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_10_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_10_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_10_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_11_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_11_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_11_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_11_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_11_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_11_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_12_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_12_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_12_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_12_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_12_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_12_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_13_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_13_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_13_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_13_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_13_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_13_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_14_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_14_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_14_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_14_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_14_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_14_6<=((others=> (others=> (others=>'0'))));
    MULTS_3_15_1<=((others=> (others=> (others=>'0'))));
    MULTS_3_15_2<=((others=> (others=> (others=>'0'))));
    MULTS_3_15_3<=((others=> (others=> (others=>'0'))));
    MULTS_3_15_4<=((others=> (others=> (others=>'0'))));
    MULTS_3_15_5<=((others=> (others=> (others=>'0'))));
    MULTS_3_15_6<=((others=> (others=> (others=>'0'))));
    EN_SUM_MULT_3<='0';

    ADD_DEPTH_1<=((others=> (others=> (others=>'0'))));Enable_STAGE_1<='0';
    ADD_DEPTH_2<=((others=> (others=> (others=>'0'))));Enable_STAGE_2<='0';
    ADD_DEPTH_3<=((others=> (others=> (others=>'0'))));Enable_STAGE_3<='0';
    ADD_DEPTH_4<=((others=> (others=> (others=>'0'))));Enable_STAGE_4<='0';
    ADD_DEPTH_5<=((others=> (others=> (others=>'0'))));Enable_STAGE_5<='0';

    MULT_1_1<=((others=> (others=> (others=>'0'))));    MULT_1_2<=((others=> (others=> (others=>'0'))));    MULT_1_3<=((others=> (others=> (others=>'0'))));    MULT_1_4<=((others=> (others=> (others=>'0'))));    MULT_1_5<=((others=> (others=> (others=>'0'))));    MULT_1_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_1_3<=(others => '0');BIAS_1<=(others => '0');ReLU_1<=(others => '0');
    MULT_2_1<=((others=> (others=> (others=>'0'))));    MULT_2_2<=((others=> (others=> (others=>'0'))));    MULT_2_3<=((others=> (others=> (others=>'0'))));    MULT_2_4<=((others=> (others=> (others=>'0'))));    MULT_2_5<=((others=> (others=> (others=>'0'))));    MULT_2_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_2_3<=(others => '0');BIAS_2<=(others => '0');ReLU_2<=(others => '0');
    MULT_3_1<=((others=> (others=> (others=>'0'))));    MULT_3_2<=((others=> (others=> (others=>'0'))));    MULT_3_3<=((others=> (others=> (others=>'0'))));    MULT_3_4<=((others=> (others=> (others=>'0'))));    MULT_3_5<=((others=> (others=> (others=>'0'))));    MULT_3_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_3_3<=(others => '0');BIAS_3<=(others => '0');ReLU_3<=(others => '0');
    MULT_4_1<=((others=> (others=> (others=>'0'))));    MULT_4_2<=((others=> (others=> (others=>'0'))));    MULT_4_3<=((others=> (others=> (others=>'0'))));    MULT_4_4<=((others=> (others=> (others=>'0'))));    MULT_4_5<=((others=> (others=> (others=>'0'))));    MULT_4_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_4_3<=(others => '0');BIAS_4<=(others => '0');ReLU_4<=(others => '0');
    MULT_5_1<=((others=> (others=> (others=>'0'))));    MULT_5_2<=((others=> (others=> (others=>'0'))));    MULT_5_3<=((others=> (others=> (others=>'0'))));    MULT_5_4<=((others=> (others=> (others=>'0'))));    MULT_5_5<=((others=> (others=> (others=>'0'))));    MULT_5_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_5_3<=(others => '0');BIAS_5<=(others => '0');ReLU_5<=(others => '0');
    MULT_6_1<=((others=> (others=> (others=>'0'))));    MULT_6_2<=((others=> (others=> (others=>'0'))));    MULT_6_3<=((others=> (others=> (others=>'0'))));    MULT_6_4<=((others=> (others=> (others=>'0'))));    MULT_6_5<=((others=> (others=> (others=>'0'))));    MULT_6_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_6_3<=(others => '0');BIAS_6<=(others => '0');ReLU_6<=(others => '0');
    MULT_7_1<=((others=> (others=> (others=>'0'))));    MULT_7_2<=((others=> (others=> (others=>'0'))));    MULT_7_3<=((others=> (others=> (others=>'0'))));    MULT_7_4<=((others=> (others=> (others=>'0'))));    MULT_7_5<=((others=> (others=> (others=>'0'))));    MULT_7_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_7_3<=(others => '0');BIAS_7<=(others => '0');ReLU_7<=(others => '0');
    MULT_8_1<=((others=> (others=> (others=>'0'))));    MULT_8_2<=((others=> (others=> (others=>'0'))));    MULT_8_3<=((others=> (others=> (others=>'0'))));    MULT_8_4<=((others=> (others=> (others=>'0'))));    MULT_8_5<=((others=> (others=> (others=>'0'))));    MULT_8_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_8_3<=(others => '0');BIAS_8<=(others => '0');ReLU_8<=(others => '0');
    MULT_9_1<=((others=> (others=> (others=>'0'))));    MULT_9_2<=((others=> (others=> (others=>'0'))));    MULT_9_3<=((others=> (others=> (others=>'0'))));    MULT_9_4<=((others=> (others=> (others=>'0'))));    MULT_9_5<=((others=> (others=> (others=>'0'))));    MULT_9_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_9_3<=(others => '0');BIAS_9<=(others => '0');ReLU_9<=(others => '0');
    MULT_10_1<=((others=> (others=> (others=>'0'))));    MULT_10_2<=((others=> (others=> (others=>'0'))));    MULT_10_3<=((others=> (others=> (others=>'0'))));    MULT_10_4<=((others=> (others=> (others=>'0'))));    MULT_10_5<=((others=> (others=> (others=>'0'))));    MULT_10_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_10_3<=(others => '0');BIAS_10<=(others => '0');ReLU_10<=(others => '0');
    MULT_11_1<=((others=> (others=> (others=>'0'))));    MULT_11_2<=((others=> (others=> (others=>'0'))));    MULT_11_3<=((others=> (others=> (others=>'0'))));    MULT_11_4<=((others=> (others=> (others=>'0'))));    MULT_11_5<=((others=> (others=> (others=>'0'))));    MULT_11_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_11_3<=(others => '0');BIAS_11<=(others => '0');ReLU_11<=(others => '0');
    MULT_12_1<=((others=> (others=> (others=>'0'))));    MULT_12_2<=((others=> (others=> (others=>'0'))));    MULT_12_3<=((others=> (others=> (others=>'0'))));    MULT_12_4<=((others=> (others=> (others=>'0'))));    MULT_12_5<=((others=> (others=> (others=>'0'))));    MULT_12_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_12_3<=(others => '0');BIAS_12<=(others => '0');ReLU_12<=(others => '0');
    MULT_13_1<=((others=> (others=> (others=>'0'))));    MULT_13_2<=((others=> (others=> (others=>'0'))));    MULT_13_3<=((others=> (others=> (others=>'0'))));    MULT_13_4<=((others=> (others=> (others=>'0'))));    MULT_13_5<=((others=> (others=> (others=>'0'))));    MULT_13_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_13_3<=(others => '0');BIAS_13<=(others => '0');ReLU_13<=(others => '0');
    MULT_14_1<=((others=> (others=> (others=>'0'))));    MULT_14_2<=((others=> (others=> (others=>'0'))));    MULT_14_3<=((others=> (others=> (others=>'0'))));    MULT_14_4<=((others=> (others=> (others=>'0'))));    MULT_14_5<=((others=> (others=> (others=>'0'))));    MULT_14_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_14_3<=(others => '0');BIAS_14<=(others => '0');ReLU_14<=(others => '0');
    MULT_15_1<=((others=> (others=> (others=>'0'))));    MULT_15_2<=((others=> (others=> (others=>'0'))));    MULT_15_3<=((others=> (others=> (others=>'0'))));    MULT_15_4<=((others=> (others=> (others=>'0'))));    MULT_15_5<=((others=> (others=> (others=>'0'))));    MULT_15_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_15_3<=(others => '0');BIAS_15<=(others => '0');ReLU_15<=(others => '0');
    MULT_16_1<=((others=> (others=> (others=>'0'))));    MULT_16_2<=((others=> (others=> (others=>'0'))));    MULT_16_3<=((others=> (others=> (others=>'0'))));    MULT_16_4<=((others=> (others=> (others=>'0'))));    MULT_16_5<=((others=> (others=> (others=>'0'))));    MULT_16_6<=((others=> (others=> (others=>'0'))));
    DOUT_BUF_16_3<=(others => '0');BIAS_16<=(others => '0');ReLU_16<=(others => '0');

----------------- FIFO_1_1 RESET---------------
    FIFO_1_ROW_1<= ((others=> (others=>'0')));HEAD_1_1<=0;TAIL_1_1<=0;
    WriteEn_1_1<= '0';ReadEn_1_1<= '0';Async_Mode_1_1<= false;
----------------- FIFO_1_2 RESET---------------
    FIFO_1_ROW_2<= ((others=> (others=>'0')));HEAD_1_2<=0;TAIL_1_2<=0;
    WriteEn_1_2<= '0';ReadEn_1_2<= '0';Async_Mode_1_2<= false;
----------------- FIFO_1_3 RESET---------------
    FIFO_1_ROW_3<= ((others=> (others=>'0')));HEAD_1_3<=0;TAIL_1_3<=0;
    WriteEn_1_3<= '0';ReadEn_1_3<= '0';Async_Mode_1_3<= false;
----------------- FIFO_1_4 RESET---------------
    FIFO_1_ROW_4<= ((others=> (others=>'0')));HEAD_1_4<=0;TAIL_1_4<=0;
    WriteEn_1_4<= '0';ReadEn_1_4<= '0';Async_Mode_1_4<= false;

----------------- FIFO_2_1 RESET---------------
    FIFO_2_ROW_1<= ((others=> (others=>'0')));HEAD_2_1<=0;TAIL_2_1<=0;
    WriteEn_2_1<= '0';ReadEn_2_1<= '0';Async_Mode_2_1<= false;
----------------- FIFO_2_2 RESET---------------
    FIFO_2_ROW_2<= ((others=> (others=>'0')));HEAD_2_2<=0;TAIL_2_2<=0;
    WriteEn_2_2<= '0';ReadEn_2_2<= '0';Async_Mode_2_2<= false;
----------------- FIFO_2_3 RESET---------------
    FIFO_2_ROW_3<= ((others=> (others=>'0')));HEAD_2_3<=0;TAIL_2_3<=0;
    WriteEn_2_3<= '0';ReadEn_2_3<= '0';Async_Mode_2_3<= false;
----------------- FIFO_2_4 RESET---------------
    FIFO_2_ROW_4<= ((others=> (others=>'0')));HEAD_2_4<=0;TAIL_2_4<=0;
    WriteEn_2_4<= '0';ReadEn_2_4<= '0';Async_Mode_2_4<= false;

----------------- FIFO_3_1 RESET---------------
    FIFO_3_ROW_1<= ((others=> (others=>'0')));HEAD_3_1<=0;TAIL_3_1<=0;
    WriteEn_3_1<= '0';ReadEn_3_1<= '0';Async_Mode_3_1<= false;
----------------- FIFO_3_2 RESET---------------
    FIFO_3_ROW_2<= ((others=> (others=>'0')));HEAD_3_2<=0;TAIL_3_2<=0;
    WriteEn_3_2<= '0';ReadEn_3_2<= '0';Async_Mode_3_2<= false;
----------------- FIFO_3_3 RESET---------------
    FIFO_3_ROW_3<= ((others=> (others=>'0')));HEAD_3_3<=0;TAIL_3_3<=0;
    WriteEn_3_3<= '0';ReadEn_3_3<= '0';Async_Mode_3_3<= false;
----------------- FIFO_3_4 RESET---------------
    FIFO_3_ROW_4<= ((others=> (others=>'0')));HEAD_3_4<=0;TAIL_3_4<=0;
    WriteEn_3_4<= '0';ReadEn_3_4<= '0';Async_Mode_3_4<= false;

----------------- FIFO_4_1 RESET---------------
    FIFO_4_ROW_1<= ((others=> (others=>'0')));HEAD_4_1<=0;TAIL_4_1<=0;
    WriteEn_4_1<= '0';ReadEn_4_1<= '0';Async_Mode_4_1<= false;
----------------- FIFO_4_2 RESET---------------
    FIFO_4_ROW_2<= ((others=> (others=>'0')));HEAD_4_2<=0;TAIL_4_2<=0;
    WriteEn_4_2<= '0';ReadEn_4_2<= '0';Async_Mode_4_2<= false;
----------------- FIFO_4_3 RESET---------------
    FIFO_4_ROW_3<= ((others=> (others=>'0')));HEAD_4_3<=0;TAIL_4_3<=0;
    WriteEn_4_3<= '0';ReadEn_4_3<= '0';Async_Mode_4_3<= false;
----------------- FIFO_4_4 RESET---------------
    FIFO_4_ROW_4<= ((others=> (others=>'0')));HEAD_4_4<=0;TAIL_4_4<=0;
    WriteEn_4_4<= '0';ReadEn_4_4<= '0';Async_Mode_4_4<= false;

----------------- FIFO_5_1 RESET---------------
    FIFO_5_ROW_1<= ((others=> (others=>'0')));HEAD_5_1<=0;TAIL_5_1<=0;
    WriteEn_5_1<= '0';ReadEn_5_1<= '0';Async_Mode_5_1<= false;
----------------- FIFO_5_2 RESET---------------
    FIFO_5_ROW_2<= ((others=> (others=>'0')));HEAD_5_2<=0;TAIL_5_2<=0;
    WriteEn_5_2<= '0';ReadEn_5_2<= '0';Async_Mode_5_2<= false;
----------------- FIFO_5_3 RESET---------------
    FIFO_5_ROW_3<= ((others=> (others=>'0')));HEAD_5_3<=0;TAIL_5_3<=0;
    WriteEn_5_3<= '0';ReadEn_5_3<= '0';Async_Mode_5_3<= false;
----------------- FIFO_5_4 RESET---------------
    FIFO_5_ROW_4<= ((others=> (others=>'0')));HEAD_5_4<=0;TAIL_5_4<=0;
    WriteEn_5_4<= '0';ReadEn_5_4<= '0';Async_Mode_5_4<= false;

----------------- FIFO_6_1 RESET---------------
    FIFO_6_ROW_1<= ((others=> (others=>'0')));HEAD_6_1<=0;TAIL_6_1<=0;
    WriteEn_6_1<= '0';ReadEn_6_1<= '0';Async_Mode_6_1<= false;
----------------- FIFO_6_2 RESET---------------
    FIFO_6_ROW_2<= ((others=> (others=>'0')));HEAD_6_2<=0;TAIL_6_2<=0;
    WriteEn_6_2<= '0';ReadEn_6_2<= '0';Async_Mode_6_2<= false;
----------------- FIFO_6_3 RESET---------------
    FIFO_6_ROW_3<= ((others=> (others=>'0')));HEAD_6_3<=0;TAIL_6_3<=0;
    WriteEn_6_3<= '0';ReadEn_6_3<= '0';Async_Mode_6_3<= false;
----------------- FIFO_6_4 RESET---------------
    FIFO_6_ROW_4<= ((others=> (others=>'0')));HEAD_6_4<=0;TAIL_6_4<=0;
    WriteEn_6_4<= '0';ReadEn_6_4<= '0';Async_Mode_6_4<= false;




------------------------------------------------ PROCESS START------------------------------------------------------
	  
   else 	
	if EN_LOC_STREAM_3='1' and EN_STREAM= '1' and OUT_PIXEL_COUNT<VALID_CYCLES  then    -- check valid data and enable stream
		
		if  FRST_TIM_EN_3='1' then EN_NXT_LYR_3<='1';end if;


               WINDOW_1(0,0)<=DIN_1_3;
               WINDOW_1(0,1)<=WINDOW_1(0,0);
               WINDOW_1(0,2)<=WINDOW_1(0,1);
               WINDOW_1(0,3)<=WINDOW_1(0,2);
               WINDOW_1(0,4)<=WINDOW_1(0,3);

               WINDOW_1(1,1)<=WINDOW_1(1,0);
               WINDOW_1(1,2)<=WINDOW_1(1,1);
               WINDOW_1(1,3)<=WINDOW_1(1,2);
               WINDOW_1(1,4)<=WINDOW_1(1,3);

               WINDOW_1(2,1)<=WINDOW_1(2,0);
               WINDOW_1(2,2)<=WINDOW_1(2,1);
               WINDOW_1(2,3)<=WINDOW_1(2,2);
               WINDOW_1(2,4)<=WINDOW_1(2,3);

               WINDOW_1(3,1)<=WINDOW_1(3,0);
               WINDOW_1(3,2)<=WINDOW_1(3,1);
               WINDOW_1(3,3)<=WINDOW_1(3,2);
               WINDOW_1(3,4)<=WINDOW_1(3,3);

               WINDOW_1(4,1)<=WINDOW_1(4,0);
               WINDOW_1(4,2)<=WINDOW_1(4,1);
               WINDOW_1(4,3)<=WINDOW_1(4,2);
               WINDOW_1(4,4)<=WINDOW_1(4,3);



               WINDOW_2(0,0)<=DIN_2_3;
               WINDOW_2(0,1)<=WINDOW_2(0,0);
               WINDOW_2(0,2)<=WINDOW_2(0,1);
               WINDOW_2(0,3)<=WINDOW_2(0,2);
               WINDOW_2(0,4)<=WINDOW_2(0,3);

               WINDOW_2(1,1)<=WINDOW_2(1,0);
               WINDOW_2(1,2)<=WINDOW_2(1,1);
               WINDOW_2(1,3)<=WINDOW_2(1,2);
               WINDOW_2(1,4)<=WINDOW_2(1,3);

               WINDOW_2(2,1)<=WINDOW_2(2,0);
               WINDOW_2(2,2)<=WINDOW_2(2,1);
               WINDOW_2(2,3)<=WINDOW_2(2,2);
               WINDOW_2(2,4)<=WINDOW_2(2,3);

               WINDOW_2(3,1)<=WINDOW_2(3,0);
               WINDOW_2(3,2)<=WINDOW_2(3,1);
               WINDOW_2(3,3)<=WINDOW_2(3,2);
               WINDOW_2(3,4)<=WINDOW_2(3,3);

               WINDOW_2(4,1)<=WINDOW_2(4,0);
               WINDOW_2(4,2)<=WINDOW_2(4,1);
               WINDOW_2(4,3)<=WINDOW_2(4,2);
               WINDOW_2(4,4)<=WINDOW_2(4,3);



               WINDOW_3(0,0)<=DIN_3_3;
               WINDOW_3(0,1)<=WINDOW_3(0,0);
               WINDOW_3(0,2)<=WINDOW_3(0,1);
               WINDOW_3(0,3)<=WINDOW_3(0,2);
               WINDOW_3(0,4)<=WINDOW_3(0,3);

               WINDOW_3(1,1)<=WINDOW_3(1,0);
               WINDOW_3(1,2)<=WINDOW_3(1,1);
               WINDOW_3(1,3)<=WINDOW_3(1,2);
               WINDOW_3(1,4)<=WINDOW_3(1,3);

               WINDOW_3(2,1)<=WINDOW_3(2,0);
               WINDOW_3(2,2)<=WINDOW_3(2,1);
               WINDOW_3(2,3)<=WINDOW_3(2,2);
               WINDOW_3(2,4)<=WINDOW_3(2,3);

               WINDOW_3(3,1)<=WINDOW_3(3,0);
               WINDOW_3(3,2)<=WINDOW_3(3,1);
               WINDOW_3(3,3)<=WINDOW_3(3,2);
               WINDOW_3(3,4)<=WINDOW_3(3,3);

               WINDOW_3(4,1)<=WINDOW_3(4,0);
               WINDOW_3(4,2)<=WINDOW_3(4,1);
               WINDOW_3(4,3)<=WINDOW_3(4,2);
               WINDOW_3(4,4)<=WINDOW_3(4,3);



               WINDOW_4(0,0)<=DIN_4_3;
               WINDOW_4(0,1)<=WINDOW_4(0,0);
               WINDOW_4(0,2)<=WINDOW_4(0,1);
               WINDOW_4(0,3)<=WINDOW_4(0,2);
               WINDOW_4(0,4)<=WINDOW_4(0,3);

               WINDOW_4(1,1)<=WINDOW_4(1,0);
               WINDOW_4(1,2)<=WINDOW_4(1,1);
               WINDOW_4(1,3)<=WINDOW_4(1,2);
               WINDOW_4(1,4)<=WINDOW_4(1,3);

               WINDOW_4(2,1)<=WINDOW_4(2,0);
               WINDOW_4(2,2)<=WINDOW_4(2,1);
               WINDOW_4(2,3)<=WINDOW_4(2,2);
               WINDOW_4(2,4)<=WINDOW_4(2,3);

               WINDOW_4(3,1)<=WINDOW_4(3,0);
               WINDOW_4(3,2)<=WINDOW_4(3,1);
               WINDOW_4(3,3)<=WINDOW_4(3,2);
               WINDOW_4(3,4)<=WINDOW_4(3,3);

               WINDOW_4(4,1)<=WINDOW_4(4,0);
               WINDOW_4(4,2)<=WINDOW_4(4,1);
               WINDOW_4(4,3)<=WINDOW_4(4,2);
               WINDOW_4(4,4)<=WINDOW_4(4,3);



               WINDOW_5(0,0)<=DIN_5_3;
               WINDOW_5(0,1)<=WINDOW_5(0,0);
               WINDOW_5(0,2)<=WINDOW_5(0,1);
               WINDOW_5(0,3)<=WINDOW_5(0,2);
               WINDOW_5(0,4)<=WINDOW_5(0,3);

               WINDOW_5(1,1)<=WINDOW_5(1,0);
               WINDOW_5(1,2)<=WINDOW_5(1,1);
               WINDOW_5(1,3)<=WINDOW_5(1,2);
               WINDOW_5(1,4)<=WINDOW_5(1,3);

               WINDOW_5(2,1)<=WINDOW_5(2,0);
               WINDOW_5(2,2)<=WINDOW_5(2,1);
               WINDOW_5(2,3)<=WINDOW_5(2,2);
               WINDOW_5(2,4)<=WINDOW_5(2,3);

               WINDOW_5(3,1)<=WINDOW_5(3,0);
               WINDOW_5(3,2)<=WINDOW_5(3,1);
               WINDOW_5(3,3)<=WINDOW_5(3,2);
               WINDOW_5(3,4)<=WINDOW_5(3,3);

               WINDOW_5(4,1)<=WINDOW_5(4,0);
               WINDOW_5(4,2)<=WINDOW_5(4,1);
               WINDOW_5(4,3)<=WINDOW_5(4,2);
               WINDOW_5(4,4)<=WINDOW_5(4,3);



               WINDOW_6(0,0)<=DIN_6_3;
               WINDOW_6(0,1)<=WINDOW_6(0,0);
               WINDOW_6(0,2)<=WINDOW_6(0,1);
               WINDOW_6(0,3)<=WINDOW_6(0,2);
               WINDOW_6(0,4)<=WINDOW_6(0,3);

               WINDOW_6(1,1)<=WINDOW_6(1,0);
               WINDOW_6(1,2)<=WINDOW_6(1,1);
               WINDOW_6(1,3)<=WINDOW_6(1,2);
               WINDOW_6(1,4)<=WINDOW_6(1,3);

               WINDOW_6(2,1)<=WINDOW_6(2,0);
               WINDOW_6(2,2)<=WINDOW_6(2,1);
               WINDOW_6(2,3)<=WINDOW_6(2,2);
               WINDOW_6(2,4)<=WINDOW_6(2,3);

               WINDOW_6(3,1)<=WINDOW_6(3,0);
               WINDOW_6(3,2)<=WINDOW_6(3,1);
               WINDOW_6(3,3)<=WINDOW_6(3,2);
               WINDOW_6(3,4)<=WINDOW_6(3,3);

               WINDOW_6(4,1)<=WINDOW_6(4,0);
               WINDOW_6(4,2)<=WINDOW_6(4,1);
               WINDOW_6(4,3)<=WINDOW_6(4,2);
               WINDOW_6(4,4)<=WINDOW_6(4,3);


                if PIXEL_COUNT=(F_SIZE-1) then
                WriteEn_1_1 <= '1';
                WriteEn_2_1 <= '1';
                WriteEn_3_1 <= '1';
                WriteEn_4_1 <= '1';
                WriteEn_5_1 <= '1';
                WriteEn_6_1 <= '1';
                else
                PIXEL_COUNT<=PIXEL_COUNT+1;
                end if;

           ----------------- Enable Read FIFO-1-1 START -------------------
				if (ReadEn_1_1 = '1') then 
				 	  WINDOW_1(1,0) <= FIFO_1_ROW_1(TAIL_1_1);
				if(TAIL_1_1 = FIFO_DEPTH-1) then
				   	TAIL_1_1<=0;  -- Rest Tail
				elsif (TAIL_1_1 = F_SIZE-1) then WriteEn_1_2<='1'; TAIL_1_1<=TAIL_1_1+1;
				else
				  	 TAIL_1_1<=TAIL_1_1+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_1_1 END -------------------

			----------------- Enable Write to FIFO_1_1 START --------------	
				if (WriteEn_1_1 = '1') then
					FIFO_1_ROW_1(HEAD_1_1)<= WINDOW_1(0,4);
				if (HEAD_1_1 = FIFO_DEPTH - 2 and Async_Mode_1_1 = false) then				 
					ReadEn_1_1<='1';
					HEAD_1_1 <= HEAD_1_1 + 1;
					Async_Mode_1_1<= true;
				else if (HEAD_1_1 = FIFO_DEPTH -1) then
					HEAD_1_1<=0;  -- Rest Head
				else
					HEAD_1_1 <= HEAD_1_1 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_1-1 END --------------


	           ----------------- Enable Read FIFO-1-2 START -------------------
				if (ReadEn_1_2 = '1') then 
				 	  WINDOW_1(2,0) <= FIFO_1_ROW_2(TAIL_1_2);
				if(TAIL_1_2 = FIFO_DEPTH-1) then
				   	TAIL_1_2<=0;  -- Rest Tail
				elsif (TAIL_1_2 = F_SIZE-1) then WriteEn_1_3<='1'; TAIL_1_2<=TAIL_1_2+1;
				else
				  	 TAIL_1_2<=TAIL_1_2+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_1_2 END -------------------

			----------------- Enable Write to FIFO_1_2 START --------------	
				if (WriteEn_1_2 = '1') then
					FIFO_1_ROW_2(HEAD_1_2)<= WINDOW_1(1,4);
				if (HEAD_1_2 = FIFO_DEPTH - 2 and Async_Mode_1_2 = false) then				 
					ReadEn_1_2<='1';
					HEAD_1_2 <= HEAD_1_2 + 1;
					Async_Mode_1_2<= true;
				else if (HEAD_1_2 = FIFO_DEPTH -1) then
					HEAD_1_2<=0;  -- Rest Head
				else
					HEAD_1_2 <= HEAD_1_2 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_1-2 END --------------


	           ----------------- Enable Read FIFO-1-3 START -------------------
				if (ReadEn_1_3 = '1') then 
				 	  WINDOW_1(3,0) <= FIFO_1_ROW_3(TAIL_1_3);
				if(TAIL_1_3 = FIFO_DEPTH-1) then
				   	TAIL_1_3<=0;  -- Rest Tail
				elsif (TAIL_1_3 = F_SIZE-1) then WriteEn_1_4<='1'; TAIL_1_3<=TAIL_1_3+1;
				else
				  	 TAIL_1_3<=TAIL_1_3+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_1_3 END -------------------

			----------------- Enable Write to FIFO_1_3 START --------------	
				if (WriteEn_1_3 = '1') then
					FIFO_1_ROW_3(HEAD_1_3)<= WINDOW_1(2,4);
				if (HEAD_1_3 = FIFO_DEPTH - 2 and Async_Mode_1_3 = false) then				 
					ReadEn_1_3<='1';
					HEAD_1_3 <= HEAD_1_3 + 1;
					Async_Mode_1_3<= true;
				else if (HEAD_1_3 = FIFO_DEPTH -1) then
					HEAD_1_3<=0;  -- Rest Head
				else
					HEAD_1_3 <= HEAD_1_3 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_1-3 END --------------


	           ----------------- Enable Read FIFO-1-4 START -------------------
				if (ReadEn_1_4 = '1') then 
				 	  WINDOW_1(4,0) <= FIFO_1_ROW_4(TAIL_1_4);
				if(TAIL_1_4 = FIFO_DEPTH-1) then
				   	TAIL_1_4<=0;  -- Rest Tail
				elsif (TAIL_1_4 = F_SIZE-1) then Enable_MULT<='1'; TAIL_1_4<=TAIL_1_4+1;
				else
				  	 TAIL_1_4<=TAIL_1_4+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_1_4 END -------------------

			----------------- Enable Write to FIFO_1_4 START --------------	
				if (WriteEn_1_4 = '1') then
					FIFO_1_ROW_4(HEAD_1_4)<= WINDOW_1(3,4);
				if (HEAD_1_4 = FIFO_DEPTH - 2 and Async_Mode_1_4 = false) then				 
					ReadEn_1_4<='1';
					HEAD_1_4 <= HEAD_1_4 + 1;
					Async_Mode_1_4<= true;
				else if (HEAD_1_4 = FIFO_DEPTH -1) then
					HEAD_1_4<=0;  -- Rest Head
				else
					HEAD_1_4 <= HEAD_1_4 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_1-4 END --------------


	

           ----------------- Enable Read FIFO-2-1 START -------------------
				if (ReadEn_2_1 = '1') then 
				 	  WINDOW_2(1,0) <= FIFO_2_ROW_1(TAIL_2_1);
				if(TAIL_2_1 = FIFO_DEPTH-1) then
				   	TAIL_2_1<=0;  -- Rest Tail
				elsif (TAIL_2_1 = F_SIZE-1) then WriteEn_2_2<='1'; TAIL_2_1<=TAIL_2_1+1;
				else
				  	 TAIL_2_1<=TAIL_2_1+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_2_1 END -------------------

			----------------- Enable Write to FIFO_2_1 START --------------	
				if (WriteEn_2_1 = '1') then
					FIFO_2_ROW_1(HEAD_2_1)<= WINDOW_2(0,4);
				if (HEAD_2_1 = FIFO_DEPTH - 2 and Async_Mode_2_1 = false) then				 
					ReadEn_2_1<='1';
					HEAD_2_1 <= HEAD_2_1 + 1;
					Async_Mode_2_1<= true;
				else if (HEAD_2_1 = FIFO_DEPTH -1) then
					HEAD_2_1<=0;  -- Rest Head
				else
					HEAD_2_1 <= HEAD_2_1 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_2-1 END --------------


	           ----------------- Enable Read FIFO-2-2 START -------------------
				if (ReadEn_2_2 = '1') then 
				 	  WINDOW_2(2,0) <= FIFO_2_ROW_2(TAIL_2_2);
				if(TAIL_2_2 = FIFO_DEPTH-1) then
				   	TAIL_2_2<=0;  -- Rest Tail
				elsif (TAIL_2_2 = F_SIZE-1) then WriteEn_2_3<='1'; TAIL_2_2<=TAIL_2_2+1;
				else
				  	 TAIL_2_2<=TAIL_2_2+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_2_2 END -------------------

			----------------- Enable Write to FIFO_2_2 START --------------	
				if (WriteEn_2_2 = '1') then
					FIFO_2_ROW_2(HEAD_2_2)<= WINDOW_2(1,4);
				if (HEAD_2_2 = FIFO_DEPTH - 2 and Async_Mode_2_2 = false) then				 
					ReadEn_2_2<='1';
					HEAD_2_2 <= HEAD_2_2 + 1;
					Async_Mode_2_2<= true;
				else if (HEAD_2_2 = FIFO_DEPTH -1) then
					HEAD_2_2<=0;  -- Rest Head
				else
					HEAD_2_2 <= HEAD_2_2 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_2-2 END --------------


	           ----------------- Enable Read FIFO-2-3 START -------------------
				if (ReadEn_2_3 = '1') then 
				 	  WINDOW_2(3,0) <= FIFO_2_ROW_3(TAIL_2_3);
				if(TAIL_2_3 = FIFO_DEPTH-1) then
				   	TAIL_2_3<=0;  -- Rest Tail
				elsif (TAIL_2_3 = F_SIZE-1) then WriteEn_2_4<='1'; TAIL_2_3<=TAIL_2_3+1;
				else
				  	 TAIL_2_3<=TAIL_2_3+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_2_3 END -------------------

			----------------- Enable Write to FIFO_2_3 START --------------	
				if (WriteEn_2_3 = '1') then
					FIFO_2_ROW_3(HEAD_2_3)<= WINDOW_2(2,4);
				if (HEAD_2_3 = FIFO_DEPTH - 2 and Async_Mode_2_3 = false) then				 
					ReadEn_2_3<='1';
					HEAD_2_3 <= HEAD_2_3 + 1;
					Async_Mode_2_3<= true;
				else if (HEAD_2_3 = FIFO_DEPTH -1) then
					HEAD_2_3<=0;  -- Rest Head
				else
					HEAD_2_3 <= HEAD_2_3 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_2-3 END --------------


	           ----------------- Enable Read FIFO-2-4 START -------------------
				if (ReadEn_2_4 = '1') then 
				 	  WINDOW_2(4,0) <= FIFO_2_ROW_4(TAIL_2_4);
				if(TAIL_2_4 = FIFO_DEPTH-1) then
				   	TAIL_2_4<=0;  -- Rest Tail
				elsif (TAIL_2_4 = F_SIZE-1) then Enable_MULT<='1'; TAIL_2_4<=TAIL_2_4+1;
				else
				  	 TAIL_2_4<=TAIL_2_4+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_2_4 END -------------------

			----------------- Enable Write to FIFO_2_4 START --------------	
				if (WriteEn_2_4 = '1') then
					FIFO_2_ROW_4(HEAD_2_4)<= WINDOW_2(3,4);
				if (HEAD_2_4 = FIFO_DEPTH - 2 and Async_Mode_2_4 = false) then				 
					ReadEn_2_4<='1';
					HEAD_2_4 <= HEAD_2_4 + 1;
					Async_Mode_2_4<= true;
				else if (HEAD_2_4 = FIFO_DEPTH -1) then
					HEAD_2_4<=0;  -- Rest Head
				else
					HEAD_2_4 <= HEAD_2_4 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_2-4 END --------------


	

           ----------------- Enable Read FIFO-3-1 START -------------------
				if (ReadEn_3_1 = '1') then 
				 	  WINDOW_3(1,0) <= FIFO_3_ROW_1(TAIL_3_1);
				if(TAIL_3_1 = FIFO_DEPTH-1) then
				   	TAIL_3_1<=0;  -- Rest Tail
				elsif (TAIL_3_1 = F_SIZE-1) then WriteEn_3_2<='1'; TAIL_3_1<=TAIL_3_1+1;
				else
				  	 TAIL_3_1<=TAIL_3_1+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_3_1 END -------------------

			----------------- Enable Write to FIFO_3_1 START --------------	
				if (WriteEn_3_1 = '1') then
					FIFO_3_ROW_1(HEAD_3_1)<= WINDOW_3(0,4);
				if (HEAD_3_1 = FIFO_DEPTH - 2 and Async_Mode_3_1 = false) then				 
					ReadEn_3_1<='1';
					HEAD_3_1 <= HEAD_3_1 + 1;
					Async_Mode_3_1<= true;
				else if (HEAD_3_1 = FIFO_DEPTH -1) then
					HEAD_3_1<=0;  -- Rest Head
				else
					HEAD_3_1 <= HEAD_3_1 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_3-1 END --------------


	           ----------------- Enable Read FIFO-3-2 START -------------------
				if (ReadEn_3_2 = '1') then 
				 	  WINDOW_3(2,0) <= FIFO_3_ROW_2(TAIL_3_2);
				if(TAIL_3_2 = FIFO_DEPTH-1) then
				   	TAIL_3_2<=0;  -- Rest Tail
				elsif (TAIL_3_2 = F_SIZE-1) then WriteEn_3_3<='1'; TAIL_3_2<=TAIL_3_2+1;
				else
				  	 TAIL_3_2<=TAIL_3_2+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_3_2 END -------------------

			----------------- Enable Write to FIFO_3_2 START --------------	
				if (WriteEn_3_2 = '1') then
					FIFO_3_ROW_2(HEAD_3_2)<= WINDOW_3(1,4);
				if (HEAD_3_2 = FIFO_DEPTH - 2 and Async_Mode_3_2 = false) then				 
					ReadEn_3_2<='1';
					HEAD_3_2 <= HEAD_3_2 + 1;
					Async_Mode_3_2<= true;
				else if (HEAD_3_2 = FIFO_DEPTH -1) then
					HEAD_3_2<=0;  -- Rest Head
				else
					HEAD_3_2 <= HEAD_3_2 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_3-2 END --------------


	           ----------------- Enable Read FIFO-3-3 START -------------------
				if (ReadEn_3_3 = '1') then 
				 	  WINDOW_3(3,0) <= FIFO_3_ROW_3(TAIL_3_3);
				if(TAIL_3_3 = FIFO_DEPTH-1) then
				   	TAIL_3_3<=0;  -- Rest Tail
				elsif (TAIL_3_3 = F_SIZE-1) then WriteEn_3_4<='1'; TAIL_3_3<=TAIL_3_3+1;
				else
				  	 TAIL_3_3<=TAIL_3_3+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_3_3 END -------------------

			----------------- Enable Write to FIFO_3_3 START --------------	
				if (WriteEn_3_3 = '1') then
					FIFO_3_ROW_3(HEAD_3_3)<= WINDOW_3(2,4);
				if (HEAD_3_3 = FIFO_DEPTH - 2 and Async_Mode_3_3 = false) then				 
					ReadEn_3_3<='1';
					HEAD_3_3 <= HEAD_3_3 + 1;
					Async_Mode_3_3<= true;
				else if (HEAD_3_3 = FIFO_DEPTH -1) then
					HEAD_3_3<=0;  -- Rest Head
				else
					HEAD_3_3 <= HEAD_3_3 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_3-3 END --------------


	           ----------------- Enable Read FIFO-3-4 START -------------------
				if (ReadEn_3_4 = '1') then 
				 	  WINDOW_3(4,0) <= FIFO_3_ROW_4(TAIL_3_4);
				if(TAIL_3_4 = FIFO_DEPTH-1) then
				   	TAIL_3_4<=0;  -- Rest Tail
				elsif (TAIL_3_4 = F_SIZE-1) then Enable_MULT<='1'; TAIL_3_4<=TAIL_3_4+1;
				else
				  	 TAIL_3_4<=TAIL_3_4+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_3_4 END -------------------

			----------------- Enable Write to FIFO_3_4 START --------------	
				if (WriteEn_3_4 = '1') then
					FIFO_3_ROW_4(HEAD_3_4)<= WINDOW_3(3,4);
				if (HEAD_3_4 = FIFO_DEPTH - 2 and Async_Mode_3_4 = false) then				 
					ReadEn_3_4<='1';
					HEAD_3_4 <= HEAD_3_4 + 1;
					Async_Mode_3_4<= true;
				else if (HEAD_3_4 = FIFO_DEPTH -1) then
					HEAD_3_4<=0;  -- Rest Head
				else
					HEAD_3_4 <= HEAD_3_4 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_3-4 END --------------


	

           ----------------- Enable Read FIFO-4-1 START -------------------
				if (ReadEn_4_1 = '1') then 
				 	  WINDOW_4(1,0) <= FIFO_4_ROW_1(TAIL_4_1);
				if(TAIL_4_1 = FIFO_DEPTH-1) then
				   	TAIL_4_1<=0;  -- Rest Tail
				elsif (TAIL_4_1 = F_SIZE-1) then WriteEn_4_2<='1'; TAIL_4_1<=TAIL_4_1+1;
				else
				  	 TAIL_4_1<=TAIL_4_1+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_4_1 END -------------------

			----------------- Enable Write to FIFO_4_1 START --------------	
				if (WriteEn_4_1 = '1') then
					FIFO_4_ROW_1(HEAD_4_1)<= WINDOW_4(0,4);
				if (HEAD_4_1 = FIFO_DEPTH - 2 and Async_Mode_4_1 = false) then				 
					ReadEn_4_1<='1';
					HEAD_4_1 <= HEAD_4_1 + 1;
					Async_Mode_4_1<= true;
				else if (HEAD_4_1 = FIFO_DEPTH -1) then
					HEAD_4_1<=0;  -- Rest Head
				else
					HEAD_4_1 <= HEAD_4_1 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_4-1 END --------------


	           ----------------- Enable Read FIFO-4-2 START -------------------
				if (ReadEn_4_2 = '1') then 
				 	  WINDOW_4(2,0) <= FIFO_4_ROW_2(TAIL_4_2);
				if(TAIL_4_2 = FIFO_DEPTH-1) then
				   	TAIL_4_2<=0;  -- Rest Tail
				elsif (TAIL_4_2 = F_SIZE-1) then WriteEn_4_3<='1'; TAIL_4_2<=TAIL_4_2+1;
				else
				  	 TAIL_4_2<=TAIL_4_2+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_4_2 END -------------------

			----------------- Enable Write to FIFO_4_2 START --------------	
				if (WriteEn_4_2 = '1') then
					FIFO_4_ROW_2(HEAD_4_2)<= WINDOW_4(1,4);
				if (HEAD_4_2 = FIFO_DEPTH - 2 and Async_Mode_4_2 = false) then				 
					ReadEn_4_2<='1';
					HEAD_4_2 <= HEAD_4_2 + 1;
					Async_Mode_4_2<= true;
				else if (HEAD_4_2 = FIFO_DEPTH -1) then
					HEAD_4_2<=0;  -- Rest Head
				else
					HEAD_4_2 <= HEAD_4_2 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_4-2 END --------------


	           ----------------- Enable Read FIFO-4-3 START -------------------
				if (ReadEn_4_3 = '1') then 
				 	  WINDOW_4(3,0) <= FIFO_4_ROW_3(TAIL_4_3);
				if(TAIL_4_3 = FIFO_DEPTH-1) then
				   	TAIL_4_3<=0;  -- Rest Tail
				elsif (TAIL_4_3 = F_SIZE-1) then WriteEn_4_4<='1'; TAIL_4_3<=TAIL_4_3+1;
				else
				  	 TAIL_4_3<=TAIL_4_3+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_4_3 END -------------------

			----------------- Enable Write to FIFO_4_3 START --------------	
				if (WriteEn_4_3 = '1') then
					FIFO_4_ROW_3(HEAD_4_3)<= WINDOW_4(2,4);
				if (HEAD_4_3 = FIFO_DEPTH - 2 and Async_Mode_4_3 = false) then				 
					ReadEn_4_3<='1';
					HEAD_4_3 <= HEAD_4_3 + 1;
					Async_Mode_4_3<= true;
				else if (HEAD_4_3 = FIFO_DEPTH -1) then
					HEAD_4_3<=0;  -- Rest Head
				else
					HEAD_4_3 <= HEAD_4_3 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_4-3 END --------------


	           ----------------- Enable Read FIFO-4-4 START -------------------
				if (ReadEn_4_4 = '1') then 
				 	  WINDOW_4(4,0) <= FIFO_4_ROW_4(TAIL_4_4);
				if(TAIL_4_4 = FIFO_DEPTH-1) then
				   	TAIL_4_4<=0;  -- Rest Tail
				elsif (TAIL_4_4 = F_SIZE-1) then Enable_MULT<='1'; TAIL_4_4<=TAIL_4_4+1;
				else
				  	 TAIL_4_4<=TAIL_4_4+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_4_4 END -------------------

			----------------- Enable Write to FIFO_4_4 START --------------	
				if (WriteEn_4_4 = '1') then
					FIFO_4_ROW_4(HEAD_4_4)<= WINDOW_4(3,4);
				if (HEAD_4_4 = FIFO_DEPTH - 2 and Async_Mode_4_4 = false) then				 
					ReadEn_4_4<='1';
					HEAD_4_4 <= HEAD_4_4 + 1;
					Async_Mode_4_4<= true;
				else if (HEAD_4_4 = FIFO_DEPTH -1) then
					HEAD_4_4<=0;  -- Rest Head
				else
					HEAD_4_4 <= HEAD_4_4 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_4-4 END --------------


	

           ----------------- Enable Read FIFO-5-1 START -------------------
				if (ReadEn_5_1 = '1') then 
				 	  WINDOW_5(1,0) <= FIFO_5_ROW_1(TAIL_5_1);
				if(TAIL_5_1 = FIFO_DEPTH-1) then
				   	TAIL_5_1<=0;  -- Rest Tail
				elsif (TAIL_5_1 = F_SIZE-1) then WriteEn_5_2<='1'; TAIL_5_1<=TAIL_5_1+1;
				else
				  	 TAIL_5_1<=TAIL_5_1+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_5_1 END -------------------

			----------------- Enable Write to FIFO_5_1 START --------------	
				if (WriteEn_5_1 = '1') then
					FIFO_5_ROW_1(HEAD_5_1)<= WINDOW_5(0,4);
				if (HEAD_5_1 = FIFO_DEPTH - 2 and Async_Mode_5_1 = false) then				 
					ReadEn_5_1<='1';
					HEAD_5_1 <= HEAD_5_1 + 1;
					Async_Mode_5_1<= true;
				else if (HEAD_5_1 = FIFO_DEPTH -1) then
					HEAD_5_1<=0;  -- Rest Head
				else
					HEAD_5_1 <= HEAD_5_1 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_5-1 END --------------


	           ----------------- Enable Read FIFO-5-2 START -------------------
				if (ReadEn_5_2 = '1') then 
				 	  WINDOW_5(2,0) <= FIFO_5_ROW_2(TAIL_5_2);
				if(TAIL_5_2 = FIFO_DEPTH-1) then
				   	TAIL_5_2<=0;  -- Rest Tail
				elsif (TAIL_5_2 = F_SIZE-1) then WriteEn_5_3<='1'; TAIL_5_2<=TAIL_5_2+1;
				else
				  	 TAIL_5_2<=TAIL_5_2+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_5_2 END -------------------

			----------------- Enable Write to FIFO_5_2 START --------------	
				if (WriteEn_5_2 = '1') then
					FIFO_5_ROW_2(HEAD_5_2)<= WINDOW_5(1,4);
				if (HEAD_5_2 = FIFO_DEPTH - 2 and Async_Mode_5_2 = false) then				 
					ReadEn_5_2<='1';
					HEAD_5_2 <= HEAD_5_2 + 1;
					Async_Mode_5_2<= true;
				else if (HEAD_5_2 = FIFO_DEPTH -1) then
					HEAD_5_2<=0;  -- Rest Head
				else
					HEAD_5_2 <= HEAD_5_2 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_5-2 END --------------


	           ----------------- Enable Read FIFO-5-3 START -------------------
				if (ReadEn_5_3 = '1') then 
				 	  WINDOW_5(3,0) <= FIFO_5_ROW_3(TAIL_5_3);
				if(TAIL_5_3 = FIFO_DEPTH-1) then
				   	TAIL_5_3<=0;  -- Rest Tail
				elsif (TAIL_5_3 = F_SIZE-1) then WriteEn_5_4<='1'; TAIL_5_3<=TAIL_5_3+1;
				else
				  	 TAIL_5_3<=TAIL_5_3+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_5_3 END -------------------

			----------------- Enable Write to FIFO_5_3 START --------------	
				if (WriteEn_5_3 = '1') then
					FIFO_5_ROW_3(HEAD_5_3)<= WINDOW_5(2,4);
				if (HEAD_5_3 = FIFO_DEPTH - 2 and Async_Mode_5_3 = false) then				 
					ReadEn_5_3<='1';
					HEAD_5_3 <= HEAD_5_3 + 1;
					Async_Mode_5_3<= true;
				else if (HEAD_5_3 = FIFO_DEPTH -1) then
					HEAD_5_3<=0;  -- Rest Head
				else
					HEAD_5_3 <= HEAD_5_3 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_5-3 END --------------


	           ----------------- Enable Read FIFO-5-4 START -------------------
				if (ReadEn_5_4 = '1') then 
				 	  WINDOW_5(4,0) <= FIFO_5_ROW_4(TAIL_5_4);
				if(TAIL_5_4 = FIFO_DEPTH-1) then
				   	TAIL_5_4<=0;  -- Rest Tail
				elsif (TAIL_5_4 = F_SIZE-1) then Enable_MULT<='1'; TAIL_5_4<=TAIL_5_4+1;
				else
				  	 TAIL_5_4<=TAIL_5_4+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_5_4 END -------------------

			----------------- Enable Write to FIFO_5_4 START --------------	
				if (WriteEn_5_4 = '1') then
					FIFO_5_ROW_4(HEAD_5_4)<= WINDOW_5(3,4);
				if (HEAD_5_4 = FIFO_DEPTH - 2 and Async_Mode_5_4 = false) then				 
					ReadEn_5_4<='1';
					HEAD_5_4 <= HEAD_5_4 + 1;
					Async_Mode_5_4<= true;
				else if (HEAD_5_4 = FIFO_DEPTH -1) then
					HEAD_5_4<=0;  -- Rest Head
				else
					HEAD_5_4 <= HEAD_5_4 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_5-4 END --------------


	

           ----------------- Enable Read FIFO-6-1 START -------------------
				if (ReadEn_6_1 = '1') then 
				 	  WINDOW_6(1,0) <= FIFO_6_ROW_1(TAIL_6_1);
				if(TAIL_6_1 = FIFO_DEPTH-1) then
				   	TAIL_6_1<=0;  -- Rest Tail
				elsif (TAIL_6_1 = F_SIZE-1) then WriteEn_6_2<='1'; TAIL_6_1<=TAIL_6_1+1;
				else
				  	 TAIL_6_1<=TAIL_6_1+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_6_1 END -------------------

			----------------- Enable Write to FIFO_6_1 START --------------	
				if (WriteEn_6_1 = '1') then
					FIFO_6_ROW_1(HEAD_6_1)<= WINDOW_6(0,4);
				if (HEAD_6_1 = FIFO_DEPTH - 2 and Async_Mode_6_1 = false) then				 
					ReadEn_6_1<='1';
					HEAD_6_1 <= HEAD_6_1 + 1;
					Async_Mode_6_1<= true;
				else if (HEAD_6_1 = FIFO_DEPTH -1) then
					HEAD_6_1<=0;  -- Rest Head
				else
					HEAD_6_1 <= HEAD_6_1 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_6-1 END --------------


	           ----------------- Enable Read FIFO-6-2 START -------------------
				if (ReadEn_6_2 = '1') then 
				 	  WINDOW_6(2,0) <= FIFO_6_ROW_2(TAIL_6_2);
				if(TAIL_6_2 = FIFO_DEPTH-1) then
				   	TAIL_6_2<=0;  -- Rest Tail
				elsif (TAIL_6_2 = F_SIZE-1) then WriteEn_6_3<='1'; TAIL_6_2<=TAIL_6_2+1;
				else
				  	 TAIL_6_2<=TAIL_6_2+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_6_2 END -------------------

			----------------- Enable Write to FIFO_6_2 START --------------	
				if (WriteEn_6_2 = '1') then
					FIFO_6_ROW_2(HEAD_6_2)<= WINDOW_6(1,4);
				if (HEAD_6_2 = FIFO_DEPTH - 2 and Async_Mode_6_2 = false) then				 
					ReadEn_6_2<='1';
					HEAD_6_2 <= HEAD_6_2 + 1;
					Async_Mode_6_2<= true;
				else if (HEAD_6_2 = FIFO_DEPTH -1) then
					HEAD_6_2<=0;  -- Rest Head
				else
					HEAD_6_2 <= HEAD_6_2 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_6-2 END --------------


	           ----------------- Enable Read FIFO-6-3 START -------------------
				if (ReadEn_6_3 = '1') then 
				 	  WINDOW_6(3,0) <= FIFO_6_ROW_3(TAIL_6_3);
				if(TAIL_6_3 = FIFO_DEPTH-1) then
				   	TAIL_6_3<=0;  -- Rest Tail
				elsif (TAIL_6_3 = F_SIZE-1) then WriteEn_6_4<='1'; TAIL_6_3<=TAIL_6_3+1;
				else
				  	 TAIL_6_3<=TAIL_6_3+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_6_3 END -------------------

			----------------- Enable Write to FIFO_6_3 START --------------	
				if (WriteEn_6_3 = '1') then
					FIFO_6_ROW_3(HEAD_6_3)<= WINDOW_6(2,4);
				if (HEAD_6_3 = FIFO_DEPTH - 2 and Async_Mode_6_3 = false) then				 
					ReadEn_6_3<='1';
					HEAD_6_3 <= HEAD_6_3 + 1;
					Async_Mode_6_3<= true;
				else if (HEAD_6_3 = FIFO_DEPTH -1) then
					HEAD_6_3<=0;  -- Rest Head
				else
					HEAD_6_3 <= HEAD_6_3 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_6-3 END --------------


	           ----------------- Enable Read FIFO-6-4 START -------------------
				if (ReadEn_6_4 = '1') then 
				 	  WINDOW_6(4,0) <= FIFO_6_ROW_4(TAIL_6_4);
				if(TAIL_6_4 = FIFO_DEPTH-1) then
				   	TAIL_6_4<=0;  -- Rest Tail
				elsif (TAIL_6_4 = F_SIZE-1) then Enable_MULT<='1'; TAIL_6_4<=TAIL_6_4+1;
				else
				  	 TAIL_6_4<=TAIL_6_4+1;
				end if;
				end if;	
			----------------- Enable Read FIFO_6_4 END -------------------

			----------------- Enable Write to FIFO_6_4 START --------------	
				if (WriteEn_6_4 = '1') then
					FIFO_6_ROW_4(HEAD_6_4)<= WINDOW_6(3,4);
				if (HEAD_6_4 = FIFO_DEPTH - 2 and Async_Mode_6_4 = false) then				 
					ReadEn_6_4<='1';
					HEAD_6_4 <= HEAD_6_4 + 1;
					Async_Mode_6_4<= true;
				else if (HEAD_6_4 = FIFO_DEPTH -1) then
					HEAD_6_4<=0;  -- Rest Head
				else
					HEAD_6_4 <= HEAD_6_4 + 1;
				end if;
				end if;
				end if;
			----------------- Enable Write to FIFO_6-4 END --------------


	

      -------------------------------------------- Enable MULT START --------------------------------------------				
	
		if Enable_MULT='1' then
			------------------------ NAME OF MULT CORROSPONDS TO WEIGHT INDEX------------------------
			MULT_1_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_1(0,0));
			MULT_1_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_1(0,0));
			MULT_1_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_1(0,0));
			MULT_1_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_1(0,0));
			MULT_1_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_1(0,0));
			MULT_1_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_1(0,0));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_2(0,0));
			MULT_2_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_2(0,0));
			MULT_2_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_2(0,0));
			MULT_2_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_2(0,0));
			MULT_2_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_2(0,0));
			MULT_2_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_2(0,0));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_3(0,0));
			MULT_3_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_3(0,0));
			MULT_3_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_3(0,0));
			MULT_3_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_3(0,0));
			MULT_3_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_3(0,0));
			MULT_3_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_3(0,0));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_4(0,0));
			MULT_4_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_4(0,0));
			MULT_4_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_4(0,0));
			MULT_4_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_4(0,0));
			MULT_4_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_4(0,0));
			MULT_4_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_4(0,0));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_5(0,0));
			MULT_5_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_5(0,0));
			MULT_5_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_5(0,0));
			MULT_5_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_5(0,0));
			MULT_5_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_5(0,0));
			MULT_5_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_5(0,0));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_6(0,0));
			MULT_6_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_6(0,0));
			MULT_6_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_6(0,0));
			MULT_6_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_6(0,0));
			MULT_6_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_6(0,0));
			MULT_6_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_6(0,0));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_7(0,0));
			MULT_7_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_7(0,0));
			MULT_7_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_7(0,0));
			MULT_7_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_7(0,0));
			MULT_7_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_7(0,0));
			MULT_7_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_7(0,0));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_8(0,0));
			MULT_8_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_8(0,0));
			MULT_8_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_8(0,0));
			MULT_8_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_8(0,0));
			MULT_8_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_8(0,0));
			MULT_8_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_8(0,0));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_9(0,0));
			MULT_9_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_9(0,0));
			MULT_9_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_9(0,0));
			MULT_9_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_9(0,0));
			MULT_9_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_9(0,0));
			MULT_9_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_9(0,0));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_10(0,0));
			MULT_10_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_10(0,0));
			MULT_10_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_10(0,0));
			MULT_10_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_10(0,0));
			MULT_10_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_10(0,0));
			MULT_10_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_10(0,0));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_11(0,0));
			MULT_11_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_11(0,0));
			MULT_11_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_11(0,0));
			MULT_11_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_11(0,0));
			MULT_11_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_11(0,0));
			MULT_11_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_11(0,0));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_12(0,0));
			MULT_12_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_12(0,0));
			MULT_12_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_12(0,0));
			MULT_12_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_12(0,0));
			MULT_12_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_12(0,0));
			MULT_12_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_12(0,0));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_13(0,0));
			MULT_13_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_13(0,0));
			MULT_13_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_13(0,0));
			MULT_13_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_13(0,0));
			MULT_13_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_13(0,0));
			MULT_13_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_13(0,0));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_14(0,0));
			MULT_14_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_14(0,0));
			MULT_14_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_14(0,0));
			MULT_14_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_14(0,0));
			MULT_14_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_14(0,0));
			MULT_14_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_14(0,0));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_15(0,0));
			MULT_15_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_15(0,0));
			MULT_15_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_15(0,0));
			MULT_15_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_15(0,0));
			MULT_15_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_15(0,0));
			MULT_15_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_15(0,0));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(0,0)<=signed(WINDOW_1(4,4))*signed(FMAP_1_16(0,0));
			MULT_16_2(0,0)<=signed(WINDOW_2(4,4))*signed(FMAP_2_16(0,0));
			MULT_16_3(0,0)<=signed(WINDOW_3(4,4))*signed(FMAP_3_16(0,0));
			MULT_16_4(0,0)<=signed(WINDOW_4(4,4))*signed(FMAP_4_16(0,0));
			MULT_16_5(0,0)<=signed(WINDOW_5(4,4))*signed(FMAP_5_16(0,0));
			MULT_16_6(0,0)<=signed(WINDOW_6(4,4))*signed(FMAP_6_16(0,0));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(0,0) -----------------------

			MULT_1_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_1(0,1));
			MULT_1_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_1(0,1));
			MULT_1_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_1(0,1));
			MULT_1_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_1(0,1));
			MULT_1_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_1(0,1));
			MULT_1_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_1(0,1));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_2(0,1));
			MULT_2_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_2(0,1));
			MULT_2_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_2(0,1));
			MULT_2_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_2(0,1));
			MULT_2_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_2(0,1));
			MULT_2_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_2(0,1));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_3(0,1));
			MULT_3_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_3(0,1));
			MULT_3_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_3(0,1));
			MULT_3_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_3(0,1));
			MULT_3_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_3(0,1));
			MULT_3_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_3(0,1));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_4(0,1));
			MULT_4_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_4(0,1));
			MULT_4_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_4(0,1));
			MULT_4_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_4(0,1));
			MULT_4_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_4(0,1));
			MULT_4_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_4(0,1));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_5(0,1));
			MULT_5_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_5(0,1));
			MULT_5_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_5(0,1));
			MULT_5_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_5(0,1));
			MULT_5_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_5(0,1));
			MULT_5_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_5(0,1));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_6(0,1));
			MULT_6_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_6(0,1));
			MULT_6_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_6(0,1));
			MULT_6_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_6(0,1));
			MULT_6_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_6(0,1));
			MULT_6_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_6(0,1));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_7(0,1));
			MULT_7_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_7(0,1));
			MULT_7_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_7(0,1));
			MULT_7_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_7(0,1));
			MULT_7_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_7(0,1));
			MULT_7_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_7(0,1));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_8(0,1));
			MULT_8_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_8(0,1));
			MULT_8_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_8(0,1));
			MULT_8_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_8(0,1));
			MULT_8_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_8(0,1));
			MULT_8_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_8(0,1));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_9(0,1));
			MULT_9_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_9(0,1));
			MULT_9_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_9(0,1));
			MULT_9_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_9(0,1));
			MULT_9_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_9(0,1));
			MULT_9_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_9(0,1));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_10(0,1));
			MULT_10_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_10(0,1));
			MULT_10_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_10(0,1));
			MULT_10_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_10(0,1));
			MULT_10_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_10(0,1));
			MULT_10_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_10(0,1));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_11(0,1));
			MULT_11_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_11(0,1));
			MULT_11_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_11(0,1));
			MULT_11_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_11(0,1));
			MULT_11_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_11(0,1));
			MULT_11_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_11(0,1));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_12(0,1));
			MULT_12_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_12(0,1));
			MULT_12_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_12(0,1));
			MULT_12_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_12(0,1));
			MULT_12_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_12(0,1));
			MULT_12_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_12(0,1));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_13(0,1));
			MULT_13_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_13(0,1));
			MULT_13_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_13(0,1));
			MULT_13_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_13(0,1));
			MULT_13_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_13(0,1));
			MULT_13_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_13(0,1));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_14(0,1));
			MULT_14_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_14(0,1));
			MULT_14_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_14(0,1));
			MULT_14_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_14(0,1));
			MULT_14_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_14(0,1));
			MULT_14_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_14(0,1));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_15(0,1));
			MULT_15_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_15(0,1));
			MULT_15_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_15(0,1));
			MULT_15_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_15(0,1));
			MULT_15_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_15(0,1));
			MULT_15_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_15(0,1));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(0,1)<=signed(WINDOW_1(4,3))*signed(FMAP_1_16(0,1));
			MULT_16_2(0,1)<=signed(WINDOW_2(4,3))*signed(FMAP_2_16(0,1));
			MULT_16_3(0,1)<=signed(WINDOW_3(4,3))*signed(FMAP_3_16(0,1));
			MULT_16_4(0,1)<=signed(WINDOW_4(4,3))*signed(FMAP_4_16(0,1));
			MULT_16_5(0,1)<=signed(WINDOW_5(4,3))*signed(FMAP_5_16(0,1));
			MULT_16_6(0,1)<=signed(WINDOW_6(4,3))*signed(FMAP_6_16(0,1));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(0,1) -----------------------

			MULT_1_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_1(0,2));
			MULT_1_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_1(0,2));
			MULT_1_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_1(0,2));
			MULT_1_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_1(0,2));
			MULT_1_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_1(0,2));
			MULT_1_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_1(0,2));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_2(0,2));
			MULT_2_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_2(0,2));
			MULT_2_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_2(0,2));
			MULT_2_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_2(0,2));
			MULT_2_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_2(0,2));
			MULT_2_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_2(0,2));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_3(0,2));
			MULT_3_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_3(0,2));
			MULT_3_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_3(0,2));
			MULT_3_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_3(0,2));
			MULT_3_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_3(0,2));
			MULT_3_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_3(0,2));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_4(0,2));
			MULT_4_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_4(0,2));
			MULT_4_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_4(0,2));
			MULT_4_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_4(0,2));
			MULT_4_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_4(0,2));
			MULT_4_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_4(0,2));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_5(0,2));
			MULT_5_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_5(0,2));
			MULT_5_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_5(0,2));
			MULT_5_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_5(0,2));
			MULT_5_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_5(0,2));
			MULT_5_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_5(0,2));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_6(0,2));
			MULT_6_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_6(0,2));
			MULT_6_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_6(0,2));
			MULT_6_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_6(0,2));
			MULT_6_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_6(0,2));
			MULT_6_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_6(0,2));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_7(0,2));
			MULT_7_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_7(0,2));
			MULT_7_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_7(0,2));
			MULT_7_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_7(0,2));
			MULT_7_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_7(0,2));
			MULT_7_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_7(0,2));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_8(0,2));
			MULT_8_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_8(0,2));
			MULT_8_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_8(0,2));
			MULT_8_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_8(0,2));
			MULT_8_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_8(0,2));
			MULT_8_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_8(0,2));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_9(0,2));
			MULT_9_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_9(0,2));
			MULT_9_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_9(0,2));
			MULT_9_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_9(0,2));
			MULT_9_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_9(0,2));
			MULT_9_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_9(0,2));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_10(0,2));
			MULT_10_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_10(0,2));
			MULT_10_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_10(0,2));
			MULT_10_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_10(0,2));
			MULT_10_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_10(0,2));
			MULT_10_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_10(0,2));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_11(0,2));
			MULT_11_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_11(0,2));
			MULT_11_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_11(0,2));
			MULT_11_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_11(0,2));
			MULT_11_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_11(0,2));
			MULT_11_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_11(0,2));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_12(0,2));
			MULT_12_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_12(0,2));
			MULT_12_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_12(0,2));
			MULT_12_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_12(0,2));
			MULT_12_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_12(0,2));
			MULT_12_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_12(0,2));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_13(0,2));
			MULT_13_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_13(0,2));
			MULT_13_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_13(0,2));
			MULT_13_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_13(0,2));
			MULT_13_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_13(0,2));
			MULT_13_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_13(0,2));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_14(0,2));
			MULT_14_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_14(0,2));
			MULT_14_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_14(0,2));
			MULT_14_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_14(0,2));
			MULT_14_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_14(0,2));
			MULT_14_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_14(0,2));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_15(0,2));
			MULT_15_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_15(0,2));
			MULT_15_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_15(0,2));
			MULT_15_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_15(0,2));
			MULT_15_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_15(0,2));
			MULT_15_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_15(0,2));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(0,2)<=signed(WINDOW_1(4,2))*signed(FMAP_1_16(0,2));
			MULT_16_2(0,2)<=signed(WINDOW_2(4,2))*signed(FMAP_2_16(0,2));
			MULT_16_3(0,2)<=signed(WINDOW_3(4,2))*signed(FMAP_3_16(0,2));
			MULT_16_4(0,2)<=signed(WINDOW_4(4,2))*signed(FMAP_4_16(0,2));
			MULT_16_5(0,2)<=signed(WINDOW_5(4,2))*signed(FMAP_5_16(0,2));
			MULT_16_6(0,2)<=signed(WINDOW_6(4,2))*signed(FMAP_6_16(0,2));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(0,2) -----------------------

			MULT_1_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_1(0,3));
			MULT_1_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_1(0,3));
			MULT_1_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_1(0,3));
			MULT_1_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_1(0,3));
			MULT_1_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_1(0,3));
			MULT_1_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_1(0,3));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_2(0,3));
			MULT_2_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_2(0,3));
			MULT_2_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_2(0,3));
			MULT_2_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_2(0,3));
			MULT_2_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_2(0,3));
			MULT_2_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_2(0,3));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_3(0,3));
			MULT_3_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_3(0,3));
			MULT_3_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_3(0,3));
			MULT_3_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_3(0,3));
			MULT_3_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_3(0,3));
			MULT_3_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_3(0,3));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_4(0,3));
			MULT_4_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_4(0,3));
			MULT_4_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_4(0,3));
			MULT_4_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_4(0,3));
			MULT_4_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_4(0,3));
			MULT_4_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_4(0,3));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_5(0,3));
			MULT_5_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_5(0,3));
			MULT_5_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_5(0,3));
			MULT_5_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_5(0,3));
			MULT_5_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_5(0,3));
			MULT_5_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_5(0,3));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_6(0,3));
			MULT_6_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_6(0,3));
			MULT_6_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_6(0,3));
			MULT_6_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_6(0,3));
			MULT_6_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_6(0,3));
			MULT_6_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_6(0,3));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_7(0,3));
			MULT_7_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_7(0,3));
			MULT_7_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_7(0,3));
			MULT_7_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_7(0,3));
			MULT_7_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_7(0,3));
			MULT_7_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_7(0,3));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_8(0,3));
			MULT_8_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_8(0,3));
			MULT_8_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_8(0,3));
			MULT_8_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_8(0,3));
			MULT_8_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_8(0,3));
			MULT_8_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_8(0,3));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_9(0,3));
			MULT_9_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_9(0,3));
			MULT_9_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_9(0,3));
			MULT_9_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_9(0,3));
			MULT_9_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_9(0,3));
			MULT_9_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_9(0,3));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_10(0,3));
			MULT_10_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_10(0,3));
			MULT_10_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_10(0,3));
			MULT_10_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_10(0,3));
			MULT_10_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_10(0,3));
			MULT_10_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_10(0,3));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_11(0,3));
			MULT_11_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_11(0,3));
			MULT_11_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_11(0,3));
			MULT_11_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_11(0,3));
			MULT_11_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_11(0,3));
			MULT_11_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_11(0,3));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_12(0,3));
			MULT_12_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_12(0,3));
			MULT_12_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_12(0,3));
			MULT_12_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_12(0,3));
			MULT_12_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_12(0,3));
			MULT_12_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_12(0,3));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_13(0,3));
			MULT_13_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_13(0,3));
			MULT_13_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_13(0,3));
			MULT_13_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_13(0,3));
			MULT_13_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_13(0,3));
			MULT_13_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_13(0,3));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_14(0,3));
			MULT_14_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_14(0,3));
			MULT_14_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_14(0,3));
			MULT_14_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_14(0,3));
			MULT_14_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_14(0,3));
			MULT_14_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_14(0,3));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_15(0,3));
			MULT_15_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_15(0,3));
			MULT_15_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_15(0,3));
			MULT_15_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_15(0,3));
			MULT_15_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_15(0,3));
			MULT_15_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_15(0,3));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(0,3)<=signed(WINDOW_1(4,1))*signed(FMAP_1_16(0,3));
			MULT_16_2(0,3)<=signed(WINDOW_2(4,1))*signed(FMAP_2_16(0,3));
			MULT_16_3(0,3)<=signed(WINDOW_3(4,1))*signed(FMAP_3_16(0,3));
			MULT_16_4(0,3)<=signed(WINDOW_4(4,1))*signed(FMAP_4_16(0,3));
			MULT_16_5(0,3)<=signed(WINDOW_5(4,1))*signed(FMAP_5_16(0,3));
			MULT_16_6(0,3)<=signed(WINDOW_6(4,1))*signed(FMAP_6_16(0,3));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(0,3) -----------------------

			MULT_1_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_1(0,4));
			MULT_1_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_1(0,4));
			MULT_1_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_1(0,4));
			MULT_1_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_1(0,4));
			MULT_1_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_1(0,4));
			MULT_1_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_1(0,4));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_2(0,4));
			MULT_2_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_2(0,4));
			MULT_2_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_2(0,4));
			MULT_2_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_2(0,4));
			MULT_2_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_2(0,4));
			MULT_2_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_2(0,4));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_3(0,4));
			MULT_3_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_3(0,4));
			MULT_3_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_3(0,4));
			MULT_3_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_3(0,4));
			MULT_3_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_3(0,4));
			MULT_3_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_3(0,4));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_4(0,4));
			MULT_4_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_4(0,4));
			MULT_4_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_4(0,4));
			MULT_4_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_4(0,4));
			MULT_4_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_4(0,4));
			MULT_4_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_4(0,4));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_5(0,4));
			MULT_5_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_5(0,4));
			MULT_5_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_5(0,4));
			MULT_5_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_5(0,4));
			MULT_5_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_5(0,4));
			MULT_5_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_5(0,4));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_6(0,4));
			MULT_6_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_6(0,4));
			MULT_6_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_6(0,4));
			MULT_6_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_6(0,4));
			MULT_6_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_6(0,4));
			MULT_6_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_6(0,4));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_7(0,4));
			MULT_7_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_7(0,4));
			MULT_7_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_7(0,4));
			MULT_7_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_7(0,4));
			MULT_7_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_7(0,4));
			MULT_7_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_7(0,4));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_8(0,4));
			MULT_8_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_8(0,4));
			MULT_8_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_8(0,4));
			MULT_8_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_8(0,4));
			MULT_8_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_8(0,4));
			MULT_8_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_8(0,4));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_9(0,4));
			MULT_9_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_9(0,4));
			MULT_9_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_9(0,4));
			MULT_9_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_9(0,4));
			MULT_9_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_9(0,4));
			MULT_9_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_9(0,4));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_10(0,4));
			MULT_10_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_10(0,4));
			MULT_10_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_10(0,4));
			MULT_10_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_10(0,4));
			MULT_10_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_10(0,4));
			MULT_10_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_10(0,4));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_11(0,4));
			MULT_11_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_11(0,4));
			MULT_11_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_11(0,4));
			MULT_11_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_11(0,4));
			MULT_11_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_11(0,4));
			MULT_11_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_11(0,4));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_12(0,4));
			MULT_12_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_12(0,4));
			MULT_12_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_12(0,4));
			MULT_12_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_12(0,4));
			MULT_12_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_12(0,4));
			MULT_12_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_12(0,4));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_13(0,4));
			MULT_13_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_13(0,4));
			MULT_13_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_13(0,4));
			MULT_13_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_13(0,4));
			MULT_13_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_13(0,4));
			MULT_13_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_13(0,4));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_14(0,4));
			MULT_14_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_14(0,4));
			MULT_14_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_14(0,4));
			MULT_14_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_14(0,4));
			MULT_14_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_14(0,4));
			MULT_14_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_14(0,4));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_15(0,4));
			MULT_15_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_15(0,4));
			MULT_15_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_15(0,4));
			MULT_15_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_15(0,4));
			MULT_15_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_15(0,4));
			MULT_15_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_15(0,4));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(0,4)<=signed(WINDOW_1(4,0))*signed(FMAP_1_16(0,4));
			MULT_16_2(0,4)<=signed(WINDOW_2(4,0))*signed(FMAP_2_16(0,4));
			MULT_16_3(0,4)<=signed(WINDOW_3(4,0))*signed(FMAP_3_16(0,4));
			MULT_16_4(0,4)<=signed(WINDOW_4(4,0))*signed(FMAP_4_16(0,4));
			MULT_16_5(0,4)<=signed(WINDOW_5(4,0))*signed(FMAP_5_16(0,4));
			MULT_16_6(0,4)<=signed(WINDOW_6(4,0))*signed(FMAP_6_16(0,4));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(0,4) -----------------------

			MULT_1_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_1(1,0));
			MULT_1_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_1(1,0));
			MULT_1_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_1(1,0));
			MULT_1_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_1(1,0));
			MULT_1_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_1(1,0));
			MULT_1_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_1(1,0));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_2(1,0));
			MULT_2_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_2(1,0));
			MULT_2_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_2(1,0));
			MULT_2_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_2(1,0));
			MULT_2_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_2(1,0));
			MULT_2_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_2(1,0));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_3(1,0));
			MULT_3_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_3(1,0));
			MULT_3_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_3(1,0));
			MULT_3_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_3(1,0));
			MULT_3_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_3(1,0));
			MULT_3_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_3(1,0));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_4(1,0));
			MULT_4_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_4(1,0));
			MULT_4_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_4(1,0));
			MULT_4_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_4(1,0));
			MULT_4_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_4(1,0));
			MULT_4_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_4(1,0));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_5(1,0));
			MULT_5_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_5(1,0));
			MULT_5_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_5(1,0));
			MULT_5_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_5(1,0));
			MULT_5_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_5(1,0));
			MULT_5_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_5(1,0));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_6(1,0));
			MULT_6_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_6(1,0));
			MULT_6_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_6(1,0));
			MULT_6_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_6(1,0));
			MULT_6_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_6(1,0));
			MULT_6_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_6(1,0));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_7(1,0));
			MULT_7_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_7(1,0));
			MULT_7_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_7(1,0));
			MULT_7_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_7(1,0));
			MULT_7_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_7(1,0));
			MULT_7_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_7(1,0));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_8(1,0));
			MULT_8_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_8(1,0));
			MULT_8_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_8(1,0));
			MULT_8_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_8(1,0));
			MULT_8_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_8(1,0));
			MULT_8_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_8(1,0));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_9(1,0));
			MULT_9_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_9(1,0));
			MULT_9_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_9(1,0));
			MULT_9_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_9(1,0));
			MULT_9_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_9(1,0));
			MULT_9_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_9(1,0));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_10(1,0));
			MULT_10_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_10(1,0));
			MULT_10_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_10(1,0));
			MULT_10_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_10(1,0));
			MULT_10_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_10(1,0));
			MULT_10_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_10(1,0));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_11(1,0));
			MULT_11_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_11(1,0));
			MULT_11_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_11(1,0));
			MULT_11_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_11(1,0));
			MULT_11_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_11(1,0));
			MULT_11_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_11(1,0));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_12(1,0));
			MULT_12_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_12(1,0));
			MULT_12_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_12(1,0));
			MULT_12_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_12(1,0));
			MULT_12_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_12(1,0));
			MULT_12_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_12(1,0));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_13(1,0));
			MULT_13_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_13(1,0));
			MULT_13_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_13(1,0));
			MULT_13_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_13(1,0));
			MULT_13_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_13(1,0));
			MULT_13_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_13(1,0));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_14(1,0));
			MULT_14_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_14(1,0));
			MULT_14_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_14(1,0));
			MULT_14_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_14(1,0));
			MULT_14_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_14(1,0));
			MULT_14_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_14(1,0));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_15(1,0));
			MULT_15_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_15(1,0));
			MULT_15_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_15(1,0));
			MULT_15_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_15(1,0));
			MULT_15_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_15(1,0));
			MULT_15_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_15(1,0));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(1,0)<=signed(WINDOW_1(3,4))*signed(FMAP_1_16(1,0));
			MULT_16_2(1,0)<=signed(WINDOW_2(3,4))*signed(FMAP_2_16(1,0));
			MULT_16_3(1,0)<=signed(WINDOW_3(3,4))*signed(FMAP_3_16(1,0));
			MULT_16_4(1,0)<=signed(WINDOW_4(3,4))*signed(FMAP_4_16(1,0));
			MULT_16_5(1,0)<=signed(WINDOW_5(3,4))*signed(FMAP_5_16(1,0));
			MULT_16_6(1,0)<=signed(WINDOW_6(3,4))*signed(FMAP_6_16(1,0));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(1,0) -----------------------

			MULT_1_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_1(1,1));
			MULT_1_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_1(1,1));
			MULT_1_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_1(1,1));
			MULT_1_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_1(1,1));
			MULT_1_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_1(1,1));
			MULT_1_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_1(1,1));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_2(1,1));
			MULT_2_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_2(1,1));
			MULT_2_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_2(1,1));
			MULT_2_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_2(1,1));
			MULT_2_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_2(1,1));
			MULT_2_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_2(1,1));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_3(1,1));
			MULT_3_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_3(1,1));
			MULT_3_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_3(1,1));
			MULT_3_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_3(1,1));
			MULT_3_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_3(1,1));
			MULT_3_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_3(1,1));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_4(1,1));
			MULT_4_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_4(1,1));
			MULT_4_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_4(1,1));
			MULT_4_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_4(1,1));
			MULT_4_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_4(1,1));
			MULT_4_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_4(1,1));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_5(1,1));
			MULT_5_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_5(1,1));
			MULT_5_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_5(1,1));
			MULT_5_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_5(1,1));
			MULT_5_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_5(1,1));
			MULT_5_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_5(1,1));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_6(1,1));
			MULT_6_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_6(1,1));
			MULT_6_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_6(1,1));
			MULT_6_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_6(1,1));
			MULT_6_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_6(1,1));
			MULT_6_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_6(1,1));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_7(1,1));
			MULT_7_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_7(1,1));
			MULT_7_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_7(1,1));
			MULT_7_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_7(1,1));
			MULT_7_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_7(1,1));
			MULT_7_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_7(1,1));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_8(1,1));
			MULT_8_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_8(1,1));
			MULT_8_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_8(1,1));
			MULT_8_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_8(1,1));
			MULT_8_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_8(1,1));
			MULT_8_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_8(1,1));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_9(1,1));
			MULT_9_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_9(1,1));
			MULT_9_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_9(1,1));
			MULT_9_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_9(1,1));
			MULT_9_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_9(1,1));
			MULT_9_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_9(1,1));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_10(1,1));
			MULT_10_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_10(1,1));
			MULT_10_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_10(1,1));
			MULT_10_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_10(1,1));
			MULT_10_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_10(1,1));
			MULT_10_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_10(1,1));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_11(1,1));
			MULT_11_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_11(1,1));
			MULT_11_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_11(1,1));
			MULT_11_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_11(1,1));
			MULT_11_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_11(1,1));
			MULT_11_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_11(1,1));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_12(1,1));
			MULT_12_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_12(1,1));
			MULT_12_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_12(1,1));
			MULT_12_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_12(1,1));
			MULT_12_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_12(1,1));
			MULT_12_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_12(1,1));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_13(1,1));
			MULT_13_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_13(1,1));
			MULT_13_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_13(1,1));
			MULT_13_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_13(1,1));
			MULT_13_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_13(1,1));
			MULT_13_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_13(1,1));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_14(1,1));
			MULT_14_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_14(1,1));
			MULT_14_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_14(1,1));
			MULT_14_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_14(1,1));
			MULT_14_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_14(1,1));
			MULT_14_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_14(1,1));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_15(1,1));
			MULT_15_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_15(1,1));
			MULT_15_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_15(1,1));
			MULT_15_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_15(1,1));
			MULT_15_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_15(1,1));
			MULT_15_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_15(1,1));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(1,1)<=signed(WINDOW_1(3,3))*signed(FMAP_1_16(1,1));
			MULT_16_2(1,1)<=signed(WINDOW_2(3,3))*signed(FMAP_2_16(1,1));
			MULT_16_3(1,1)<=signed(WINDOW_3(3,3))*signed(FMAP_3_16(1,1));
			MULT_16_4(1,1)<=signed(WINDOW_4(3,3))*signed(FMAP_4_16(1,1));
			MULT_16_5(1,1)<=signed(WINDOW_5(3,3))*signed(FMAP_5_16(1,1));
			MULT_16_6(1,1)<=signed(WINDOW_6(3,3))*signed(FMAP_6_16(1,1));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(1,1) -----------------------

			MULT_1_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_1(1,2));
			MULT_1_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_1(1,2));
			MULT_1_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_1(1,2));
			MULT_1_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_1(1,2));
			MULT_1_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_1(1,2));
			MULT_1_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_1(1,2));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_2(1,2));
			MULT_2_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_2(1,2));
			MULT_2_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_2(1,2));
			MULT_2_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_2(1,2));
			MULT_2_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_2(1,2));
			MULT_2_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_2(1,2));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_3(1,2));
			MULT_3_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_3(1,2));
			MULT_3_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_3(1,2));
			MULT_3_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_3(1,2));
			MULT_3_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_3(1,2));
			MULT_3_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_3(1,2));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_4(1,2));
			MULT_4_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_4(1,2));
			MULT_4_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_4(1,2));
			MULT_4_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_4(1,2));
			MULT_4_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_4(1,2));
			MULT_4_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_4(1,2));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_5(1,2));
			MULT_5_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_5(1,2));
			MULT_5_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_5(1,2));
			MULT_5_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_5(1,2));
			MULT_5_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_5(1,2));
			MULT_5_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_5(1,2));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_6(1,2));
			MULT_6_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_6(1,2));
			MULT_6_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_6(1,2));
			MULT_6_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_6(1,2));
			MULT_6_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_6(1,2));
			MULT_6_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_6(1,2));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_7(1,2));
			MULT_7_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_7(1,2));
			MULT_7_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_7(1,2));
			MULT_7_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_7(1,2));
			MULT_7_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_7(1,2));
			MULT_7_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_7(1,2));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_8(1,2));
			MULT_8_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_8(1,2));
			MULT_8_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_8(1,2));
			MULT_8_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_8(1,2));
			MULT_8_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_8(1,2));
			MULT_8_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_8(1,2));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_9(1,2));
			MULT_9_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_9(1,2));
			MULT_9_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_9(1,2));
			MULT_9_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_9(1,2));
			MULT_9_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_9(1,2));
			MULT_9_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_9(1,2));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_10(1,2));
			MULT_10_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_10(1,2));
			MULT_10_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_10(1,2));
			MULT_10_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_10(1,2));
			MULT_10_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_10(1,2));
			MULT_10_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_10(1,2));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_11(1,2));
			MULT_11_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_11(1,2));
			MULT_11_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_11(1,2));
			MULT_11_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_11(1,2));
			MULT_11_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_11(1,2));
			MULT_11_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_11(1,2));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_12(1,2));
			MULT_12_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_12(1,2));
			MULT_12_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_12(1,2));
			MULT_12_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_12(1,2));
			MULT_12_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_12(1,2));
			MULT_12_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_12(1,2));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_13(1,2));
			MULT_13_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_13(1,2));
			MULT_13_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_13(1,2));
			MULT_13_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_13(1,2));
			MULT_13_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_13(1,2));
			MULT_13_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_13(1,2));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_14(1,2));
			MULT_14_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_14(1,2));
			MULT_14_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_14(1,2));
			MULT_14_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_14(1,2));
			MULT_14_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_14(1,2));
			MULT_14_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_14(1,2));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_15(1,2));
			MULT_15_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_15(1,2));
			MULT_15_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_15(1,2));
			MULT_15_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_15(1,2));
			MULT_15_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_15(1,2));
			MULT_15_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_15(1,2));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(1,2)<=signed(WINDOW_1(3,2))*signed(FMAP_1_16(1,2));
			MULT_16_2(1,2)<=signed(WINDOW_2(3,2))*signed(FMAP_2_16(1,2));
			MULT_16_3(1,2)<=signed(WINDOW_3(3,2))*signed(FMAP_3_16(1,2));
			MULT_16_4(1,2)<=signed(WINDOW_4(3,2))*signed(FMAP_4_16(1,2));
			MULT_16_5(1,2)<=signed(WINDOW_5(3,2))*signed(FMAP_5_16(1,2));
			MULT_16_6(1,2)<=signed(WINDOW_6(3,2))*signed(FMAP_6_16(1,2));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(1,2) -----------------------

			MULT_1_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_1(1,3));
			MULT_1_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_1(1,3));
			MULT_1_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_1(1,3));
			MULT_1_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_1(1,3));
			MULT_1_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_1(1,3));
			MULT_1_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_1(1,3));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_2(1,3));
			MULT_2_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_2(1,3));
			MULT_2_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_2(1,3));
			MULT_2_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_2(1,3));
			MULT_2_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_2(1,3));
			MULT_2_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_2(1,3));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_3(1,3));
			MULT_3_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_3(1,3));
			MULT_3_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_3(1,3));
			MULT_3_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_3(1,3));
			MULT_3_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_3(1,3));
			MULT_3_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_3(1,3));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_4(1,3));
			MULT_4_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_4(1,3));
			MULT_4_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_4(1,3));
			MULT_4_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_4(1,3));
			MULT_4_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_4(1,3));
			MULT_4_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_4(1,3));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_5(1,3));
			MULT_5_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_5(1,3));
			MULT_5_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_5(1,3));
			MULT_5_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_5(1,3));
			MULT_5_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_5(1,3));
			MULT_5_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_5(1,3));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_6(1,3));
			MULT_6_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_6(1,3));
			MULT_6_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_6(1,3));
			MULT_6_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_6(1,3));
			MULT_6_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_6(1,3));
			MULT_6_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_6(1,3));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_7(1,3));
			MULT_7_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_7(1,3));
			MULT_7_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_7(1,3));
			MULT_7_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_7(1,3));
			MULT_7_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_7(1,3));
			MULT_7_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_7(1,3));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_8(1,3));
			MULT_8_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_8(1,3));
			MULT_8_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_8(1,3));
			MULT_8_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_8(1,3));
			MULT_8_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_8(1,3));
			MULT_8_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_8(1,3));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_9(1,3));
			MULT_9_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_9(1,3));
			MULT_9_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_9(1,3));
			MULT_9_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_9(1,3));
			MULT_9_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_9(1,3));
			MULT_9_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_9(1,3));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_10(1,3));
			MULT_10_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_10(1,3));
			MULT_10_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_10(1,3));
			MULT_10_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_10(1,3));
			MULT_10_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_10(1,3));
			MULT_10_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_10(1,3));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_11(1,3));
			MULT_11_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_11(1,3));
			MULT_11_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_11(1,3));
			MULT_11_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_11(1,3));
			MULT_11_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_11(1,3));
			MULT_11_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_11(1,3));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_12(1,3));
			MULT_12_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_12(1,3));
			MULT_12_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_12(1,3));
			MULT_12_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_12(1,3));
			MULT_12_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_12(1,3));
			MULT_12_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_12(1,3));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_13(1,3));
			MULT_13_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_13(1,3));
			MULT_13_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_13(1,3));
			MULT_13_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_13(1,3));
			MULT_13_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_13(1,3));
			MULT_13_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_13(1,3));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_14(1,3));
			MULT_14_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_14(1,3));
			MULT_14_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_14(1,3));
			MULT_14_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_14(1,3));
			MULT_14_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_14(1,3));
			MULT_14_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_14(1,3));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_15(1,3));
			MULT_15_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_15(1,3));
			MULT_15_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_15(1,3));
			MULT_15_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_15(1,3));
			MULT_15_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_15(1,3));
			MULT_15_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_15(1,3));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(1,3)<=signed(WINDOW_1(3,1))*signed(FMAP_1_16(1,3));
			MULT_16_2(1,3)<=signed(WINDOW_2(3,1))*signed(FMAP_2_16(1,3));
			MULT_16_3(1,3)<=signed(WINDOW_3(3,1))*signed(FMAP_3_16(1,3));
			MULT_16_4(1,3)<=signed(WINDOW_4(3,1))*signed(FMAP_4_16(1,3));
			MULT_16_5(1,3)<=signed(WINDOW_5(3,1))*signed(FMAP_5_16(1,3));
			MULT_16_6(1,3)<=signed(WINDOW_6(3,1))*signed(FMAP_6_16(1,3));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(1,3) -----------------------

			MULT_1_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_1(1,4));
			MULT_1_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_1(1,4));
			MULT_1_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_1(1,4));
			MULT_1_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_1(1,4));
			MULT_1_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_1(1,4));
			MULT_1_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_1(1,4));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_2(1,4));
			MULT_2_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_2(1,4));
			MULT_2_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_2(1,4));
			MULT_2_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_2(1,4));
			MULT_2_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_2(1,4));
			MULT_2_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_2(1,4));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_3(1,4));
			MULT_3_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_3(1,4));
			MULT_3_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_3(1,4));
			MULT_3_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_3(1,4));
			MULT_3_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_3(1,4));
			MULT_3_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_3(1,4));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_4(1,4));
			MULT_4_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_4(1,4));
			MULT_4_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_4(1,4));
			MULT_4_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_4(1,4));
			MULT_4_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_4(1,4));
			MULT_4_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_4(1,4));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_5(1,4));
			MULT_5_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_5(1,4));
			MULT_5_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_5(1,4));
			MULT_5_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_5(1,4));
			MULT_5_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_5(1,4));
			MULT_5_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_5(1,4));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_6(1,4));
			MULT_6_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_6(1,4));
			MULT_6_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_6(1,4));
			MULT_6_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_6(1,4));
			MULT_6_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_6(1,4));
			MULT_6_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_6(1,4));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_7(1,4));
			MULT_7_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_7(1,4));
			MULT_7_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_7(1,4));
			MULT_7_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_7(1,4));
			MULT_7_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_7(1,4));
			MULT_7_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_7(1,4));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_8(1,4));
			MULT_8_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_8(1,4));
			MULT_8_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_8(1,4));
			MULT_8_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_8(1,4));
			MULT_8_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_8(1,4));
			MULT_8_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_8(1,4));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_9(1,4));
			MULT_9_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_9(1,4));
			MULT_9_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_9(1,4));
			MULT_9_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_9(1,4));
			MULT_9_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_9(1,4));
			MULT_9_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_9(1,4));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_10(1,4));
			MULT_10_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_10(1,4));
			MULT_10_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_10(1,4));
			MULT_10_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_10(1,4));
			MULT_10_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_10(1,4));
			MULT_10_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_10(1,4));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_11(1,4));
			MULT_11_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_11(1,4));
			MULT_11_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_11(1,4));
			MULT_11_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_11(1,4));
			MULT_11_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_11(1,4));
			MULT_11_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_11(1,4));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_12(1,4));
			MULT_12_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_12(1,4));
			MULT_12_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_12(1,4));
			MULT_12_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_12(1,4));
			MULT_12_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_12(1,4));
			MULT_12_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_12(1,4));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_13(1,4));
			MULT_13_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_13(1,4));
			MULT_13_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_13(1,4));
			MULT_13_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_13(1,4));
			MULT_13_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_13(1,4));
			MULT_13_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_13(1,4));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_14(1,4));
			MULT_14_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_14(1,4));
			MULT_14_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_14(1,4));
			MULT_14_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_14(1,4));
			MULT_14_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_14(1,4));
			MULT_14_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_14(1,4));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_15(1,4));
			MULT_15_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_15(1,4));
			MULT_15_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_15(1,4));
			MULT_15_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_15(1,4));
			MULT_15_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_15(1,4));
			MULT_15_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_15(1,4));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(1,4)<=signed(WINDOW_1(3,0))*signed(FMAP_1_16(1,4));
			MULT_16_2(1,4)<=signed(WINDOW_2(3,0))*signed(FMAP_2_16(1,4));
			MULT_16_3(1,4)<=signed(WINDOW_3(3,0))*signed(FMAP_3_16(1,4));
			MULT_16_4(1,4)<=signed(WINDOW_4(3,0))*signed(FMAP_4_16(1,4));
			MULT_16_5(1,4)<=signed(WINDOW_5(3,0))*signed(FMAP_5_16(1,4));
			MULT_16_6(1,4)<=signed(WINDOW_6(3,0))*signed(FMAP_6_16(1,4));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(1,4) -----------------------

			MULT_1_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_1(2,0));
			MULT_1_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_1(2,0));
			MULT_1_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_1(2,0));
			MULT_1_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_1(2,0));
			MULT_1_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_1(2,0));
			MULT_1_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_1(2,0));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_2(2,0));
			MULT_2_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_2(2,0));
			MULT_2_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_2(2,0));
			MULT_2_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_2(2,0));
			MULT_2_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_2(2,0));
			MULT_2_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_2(2,0));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_3(2,0));
			MULT_3_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_3(2,0));
			MULT_3_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_3(2,0));
			MULT_3_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_3(2,0));
			MULT_3_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_3(2,0));
			MULT_3_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_3(2,0));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_4(2,0));
			MULT_4_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_4(2,0));
			MULT_4_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_4(2,0));
			MULT_4_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_4(2,0));
			MULT_4_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_4(2,0));
			MULT_4_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_4(2,0));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_5(2,0));
			MULT_5_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_5(2,0));
			MULT_5_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_5(2,0));
			MULT_5_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_5(2,0));
			MULT_5_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_5(2,0));
			MULT_5_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_5(2,0));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_6(2,0));
			MULT_6_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_6(2,0));
			MULT_6_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_6(2,0));
			MULT_6_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_6(2,0));
			MULT_6_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_6(2,0));
			MULT_6_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_6(2,0));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_7(2,0));
			MULT_7_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_7(2,0));
			MULT_7_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_7(2,0));
			MULT_7_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_7(2,0));
			MULT_7_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_7(2,0));
			MULT_7_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_7(2,0));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_8(2,0));
			MULT_8_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_8(2,0));
			MULT_8_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_8(2,0));
			MULT_8_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_8(2,0));
			MULT_8_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_8(2,0));
			MULT_8_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_8(2,0));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_9(2,0));
			MULT_9_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_9(2,0));
			MULT_9_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_9(2,0));
			MULT_9_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_9(2,0));
			MULT_9_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_9(2,0));
			MULT_9_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_9(2,0));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_10(2,0));
			MULT_10_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_10(2,0));
			MULT_10_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_10(2,0));
			MULT_10_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_10(2,0));
			MULT_10_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_10(2,0));
			MULT_10_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_10(2,0));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_11(2,0));
			MULT_11_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_11(2,0));
			MULT_11_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_11(2,0));
			MULT_11_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_11(2,0));
			MULT_11_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_11(2,0));
			MULT_11_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_11(2,0));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_12(2,0));
			MULT_12_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_12(2,0));
			MULT_12_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_12(2,0));
			MULT_12_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_12(2,0));
			MULT_12_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_12(2,0));
			MULT_12_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_12(2,0));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_13(2,0));
			MULT_13_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_13(2,0));
			MULT_13_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_13(2,0));
			MULT_13_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_13(2,0));
			MULT_13_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_13(2,0));
			MULT_13_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_13(2,0));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_14(2,0));
			MULT_14_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_14(2,0));
			MULT_14_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_14(2,0));
			MULT_14_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_14(2,0));
			MULT_14_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_14(2,0));
			MULT_14_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_14(2,0));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_15(2,0));
			MULT_15_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_15(2,0));
			MULT_15_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_15(2,0));
			MULT_15_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_15(2,0));
			MULT_15_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_15(2,0));
			MULT_15_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_15(2,0));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(2,0)<=signed(WINDOW_1(2,4))*signed(FMAP_1_16(2,0));
			MULT_16_2(2,0)<=signed(WINDOW_2(2,4))*signed(FMAP_2_16(2,0));
			MULT_16_3(2,0)<=signed(WINDOW_3(2,4))*signed(FMAP_3_16(2,0));
			MULT_16_4(2,0)<=signed(WINDOW_4(2,4))*signed(FMAP_4_16(2,0));
			MULT_16_5(2,0)<=signed(WINDOW_5(2,4))*signed(FMAP_5_16(2,0));
			MULT_16_6(2,0)<=signed(WINDOW_6(2,4))*signed(FMAP_6_16(2,0));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(2,0) -----------------------

			MULT_1_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_1(2,1));
			MULT_1_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_1(2,1));
			MULT_1_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_1(2,1));
			MULT_1_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_1(2,1));
			MULT_1_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_1(2,1));
			MULT_1_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_1(2,1));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_2(2,1));
			MULT_2_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_2(2,1));
			MULT_2_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_2(2,1));
			MULT_2_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_2(2,1));
			MULT_2_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_2(2,1));
			MULT_2_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_2(2,1));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_3(2,1));
			MULT_3_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_3(2,1));
			MULT_3_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_3(2,1));
			MULT_3_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_3(2,1));
			MULT_3_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_3(2,1));
			MULT_3_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_3(2,1));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_4(2,1));
			MULT_4_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_4(2,1));
			MULT_4_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_4(2,1));
			MULT_4_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_4(2,1));
			MULT_4_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_4(2,1));
			MULT_4_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_4(2,1));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_5(2,1));
			MULT_5_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_5(2,1));
			MULT_5_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_5(2,1));
			MULT_5_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_5(2,1));
			MULT_5_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_5(2,1));
			MULT_5_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_5(2,1));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_6(2,1));
			MULT_6_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_6(2,1));
			MULT_6_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_6(2,1));
			MULT_6_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_6(2,1));
			MULT_6_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_6(2,1));
			MULT_6_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_6(2,1));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_7(2,1));
			MULT_7_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_7(2,1));
			MULT_7_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_7(2,1));
			MULT_7_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_7(2,1));
			MULT_7_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_7(2,1));
			MULT_7_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_7(2,1));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_8(2,1));
			MULT_8_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_8(2,1));
			MULT_8_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_8(2,1));
			MULT_8_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_8(2,1));
			MULT_8_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_8(2,1));
			MULT_8_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_8(2,1));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_9(2,1));
			MULT_9_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_9(2,1));
			MULT_9_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_9(2,1));
			MULT_9_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_9(2,1));
			MULT_9_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_9(2,1));
			MULT_9_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_9(2,1));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_10(2,1));
			MULT_10_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_10(2,1));
			MULT_10_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_10(2,1));
			MULT_10_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_10(2,1));
			MULT_10_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_10(2,1));
			MULT_10_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_10(2,1));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_11(2,1));
			MULT_11_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_11(2,1));
			MULT_11_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_11(2,1));
			MULT_11_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_11(2,1));
			MULT_11_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_11(2,1));
			MULT_11_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_11(2,1));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_12(2,1));
			MULT_12_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_12(2,1));
			MULT_12_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_12(2,1));
			MULT_12_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_12(2,1));
			MULT_12_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_12(2,1));
			MULT_12_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_12(2,1));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_13(2,1));
			MULT_13_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_13(2,1));
			MULT_13_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_13(2,1));
			MULT_13_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_13(2,1));
			MULT_13_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_13(2,1));
			MULT_13_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_13(2,1));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_14(2,1));
			MULT_14_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_14(2,1));
			MULT_14_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_14(2,1));
			MULT_14_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_14(2,1));
			MULT_14_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_14(2,1));
			MULT_14_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_14(2,1));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_15(2,1));
			MULT_15_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_15(2,1));
			MULT_15_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_15(2,1));
			MULT_15_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_15(2,1));
			MULT_15_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_15(2,1));
			MULT_15_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_15(2,1));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(2,1)<=signed(WINDOW_1(2,3))*signed(FMAP_1_16(2,1));
			MULT_16_2(2,1)<=signed(WINDOW_2(2,3))*signed(FMAP_2_16(2,1));
			MULT_16_3(2,1)<=signed(WINDOW_3(2,3))*signed(FMAP_3_16(2,1));
			MULT_16_4(2,1)<=signed(WINDOW_4(2,3))*signed(FMAP_4_16(2,1));
			MULT_16_5(2,1)<=signed(WINDOW_5(2,3))*signed(FMAP_5_16(2,1));
			MULT_16_6(2,1)<=signed(WINDOW_6(2,3))*signed(FMAP_6_16(2,1));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(2,1) -----------------------

			MULT_1_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_1(2,2));
			MULT_1_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_1(2,2));
			MULT_1_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_1(2,2));
			MULT_1_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_1(2,2));
			MULT_1_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_1(2,2));
			MULT_1_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_1(2,2));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_2(2,2));
			MULT_2_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_2(2,2));
			MULT_2_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_2(2,2));
			MULT_2_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_2(2,2));
			MULT_2_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_2(2,2));
			MULT_2_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_2(2,2));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_3(2,2));
			MULT_3_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_3(2,2));
			MULT_3_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_3(2,2));
			MULT_3_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_3(2,2));
			MULT_3_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_3(2,2));
			MULT_3_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_3(2,2));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_4(2,2));
			MULT_4_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_4(2,2));
			MULT_4_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_4(2,2));
			MULT_4_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_4(2,2));
			MULT_4_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_4(2,2));
			MULT_4_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_4(2,2));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_5(2,2));
			MULT_5_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_5(2,2));
			MULT_5_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_5(2,2));
			MULT_5_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_5(2,2));
			MULT_5_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_5(2,2));
			MULT_5_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_5(2,2));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_6(2,2));
			MULT_6_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_6(2,2));
			MULT_6_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_6(2,2));
			MULT_6_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_6(2,2));
			MULT_6_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_6(2,2));
			MULT_6_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_6(2,2));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_7(2,2));
			MULT_7_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_7(2,2));
			MULT_7_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_7(2,2));
			MULT_7_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_7(2,2));
			MULT_7_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_7(2,2));
			MULT_7_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_7(2,2));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_8(2,2));
			MULT_8_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_8(2,2));
			MULT_8_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_8(2,2));
			MULT_8_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_8(2,2));
			MULT_8_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_8(2,2));
			MULT_8_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_8(2,2));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_9(2,2));
			MULT_9_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_9(2,2));
			MULT_9_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_9(2,2));
			MULT_9_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_9(2,2));
			MULT_9_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_9(2,2));
			MULT_9_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_9(2,2));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_10(2,2));
			MULT_10_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_10(2,2));
			MULT_10_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_10(2,2));
			MULT_10_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_10(2,2));
			MULT_10_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_10(2,2));
			MULT_10_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_10(2,2));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_11(2,2));
			MULT_11_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_11(2,2));
			MULT_11_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_11(2,2));
			MULT_11_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_11(2,2));
			MULT_11_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_11(2,2));
			MULT_11_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_11(2,2));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_12(2,2));
			MULT_12_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_12(2,2));
			MULT_12_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_12(2,2));
			MULT_12_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_12(2,2));
			MULT_12_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_12(2,2));
			MULT_12_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_12(2,2));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_13(2,2));
			MULT_13_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_13(2,2));
			MULT_13_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_13(2,2));
			MULT_13_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_13(2,2));
			MULT_13_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_13(2,2));
			MULT_13_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_13(2,2));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_14(2,2));
			MULT_14_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_14(2,2));
			MULT_14_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_14(2,2));
			MULT_14_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_14(2,2));
			MULT_14_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_14(2,2));
			MULT_14_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_14(2,2));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_15(2,2));
			MULT_15_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_15(2,2));
			MULT_15_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_15(2,2));
			MULT_15_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_15(2,2));
			MULT_15_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_15(2,2));
			MULT_15_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_15(2,2));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(2,2)<=signed(WINDOW_1(2,2))*signed(FMAP_1_16(2,2));
			MULT_16_2(2,2)<=signed(WINDOW_2(2,2))*signed(FMAP_2_16(2,2));
			MULT_16_3(2,2)<=signed(WINDOW_3(2,2))*signed(FMAP_3_16(2,2));
			MULT_16_4(2,2)<=signed(WINDOW_4(2,2))*signed(FMAP_4_16(2,2));
			MULT_16_5(2,2)<=signed(WINDOW_5(2,2))*signed(FMAP_5_16(2,2));
			MULT_16_6(2,2)<=signed(WINDOW_6(2,2))*signed(FMAP_6_16(2,2));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(2,2) -----------------------

			MULT_1_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_1(2,3));
			MULT_1_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_1(2,3));
			MULT_1_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_1(2,3));
			MULT_1_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_1(2,3));
			MULT_1_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_1(2,3));
			MULT_1_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_1(2,3));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_2(2,3));
			MULT_2_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_2(2,3));
			MULT_2_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_2(2,3));
			MULT_2_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_2(2,3));
			MULT_2_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_2(2,3));
			MULT_2_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_2(2,3));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_3(2,3));
			MULT_3_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_3(2,3));
			MULT_3_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_3(2,3));
			MULT_3_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_3(2,3));
			MULT_3_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_3(2,3));
			MULT_3_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_3(2,3));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_4(2,3));
			MULT_4_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_4(2,3));
			MULT_4_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_4(2,3));
			MULT_4_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_4(2,3));
			MULT_4_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_4(2,3));
			MULT_4_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_4(2,3));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_5(2,3));
			MULT_5_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_5(2,3));
			MULT_5_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_5(2,3));
			MULT_5_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_5(2,3));
			MULT_5_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_5(2,3));
			MULT_5_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_5(2,3));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_6(2,3));
			MULT_6_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_6(2,3));
			MULT_6_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_6(2,3));
			MULT_6_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_6(2,3));
			MULT_6_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_6(2,3));
			MULT_6_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_6(2,3));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_7(2,3));
			MULT_7_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_7(2,3));
			MULT_7_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_7(2,3));
			MULT_7_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_7(2,3));
			MULT_7_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_7(2,3));
			MULT_7_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_7(2,3));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_8(2,3));
			MULT_8_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_8(2,3));
			MULT_8_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_8(2,3));
			MULT_8_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_8(2,3));
			MULT_8_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_8(2,3));
			MULT_8_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_8(2,3));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_9(2,3));
			MULT_9_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_9(2,3));
			MULT_9_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_9(2,3));
			MULT_9_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_9(2,3));
			MULT_9_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_9(2,3));
			MULT_9_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_9(2,3));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_10(2,3));
			MULT_10_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_10(2,3));
			MULT_10_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_10(2,3));
			MULT_10_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_10(2,3));
			MULT_10_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_10(2,3));
			MULT_10_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_10(2,3));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_11(2,3));
			MULT_11_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_11(2,3));
			MULT_11_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_11(2,3));
			MULT_11_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_11(2,3));
			MULT_11_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_11(2,3));
			MULT_11_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_11(2,3));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_12(2,3));
			MULT_12_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_12(2,3));
			MULT_12_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_12(2,3));
			MULT_12_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_12(2,3));
			MULT_12_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_12(2,3));
			MULT_12_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_12(2,3));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_13(2,3));
			MULT_13_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_13(2,3));
			MULT_13_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_13(2,3));
			MULT_13_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_13(2,3));
			MULT_13_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_13(2,3));
			MULT_13_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_13(2,3));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_14(2,3));
			MULT_14_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_14(2,3));
			MULT_14_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_14(2,3));
			MULT_14_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_14(2,3));
			MULT_14_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_14(2,3));
			MULT_14_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_14(2,3));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_15(2,3));
			MULT_15_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_15(2,3));
			MULT_15_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_15(2,3));
			MULT_15_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_15(2,3));
			MULT_15_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_15(2,3));
			MULT_15_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_15(2,3));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(2,3)<=signed(WINDOW_1(2,1))*signed(FMAP_1_16(2,3));
			MULT_16_2(2,3)<=signed(WINDOW_2(2,1))*signed(FMAP_2_16(2,3));
			MULT_16_3(2,3)<=signed(WINDOW_3(2,1))*signed(FMAP_3_16(2,3));
			MULT_16_4(2,3)<=signed(WINDOW_4(2,1))*signed(FMAP_4_16(2,3));
			MULT_16_5(2,3)<=signed(WINDOW_5(2,1))*signed(FMAP_5_16(2,3));
			MULT_16_6(2,3)<=signed(WINDOW_6(2,1))*signed(FMAP_6_16(2,3));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(2,3) -----------------------

			MULT_1_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_1(2,4));
			MULT_1_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_1(2,4));
			MULT_1_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_1(2,4));
			MULT_1_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_1(2,4));
			MULT_1_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_1(2,4));
			MULT_1_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_1(2,4));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_2(2,4));
			MULT_2_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_2(2,4));
			MULT_2_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_2(2,4));
			MULT_2_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_2(2,4));
			MULT_2_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_2(2,4));
			MULT_2_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_2(2,4));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_3(2,4));
			MULT_3_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_3(2,4));
			MULT_3_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_3(2,4));
			MULT_3_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_3(2,4));
			MULT_3_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_3(2,4));
			MULT_3_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_3(2,4));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_4(2,4));
			MULT_4_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_4(2,4));
			MULT_4_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_4(2,4));
			MULT_4_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_4(2,4));
			MULT_4_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_4(2,4));
			MULT_4_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_4(2,4));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_5(2,4));
			MULT_5_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_5(2,4));
			MULT_5_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_5(2,4));
			MULT_5_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_5(2,4));
			MULT_5_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_5(2,4));
			MULT_5_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_5(2,4));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_6(2,4));
			MULT_6_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_6(2,4));
			MULT_6_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_6(2,4));
			MULT_6_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_6(2,4));
			MULT_6_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_6(2,4));
			MULT_6_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_6(2,4));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_7(2,4));
			MULT_7_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_7(2,4));
			MULT_7_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_7(2,4));
			MULT_7_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_7(2,4));
			MULT_7_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_7(2,4));
			MULT_7_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_7(2,4));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_8(2,4));
			MULT_8_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_8(2,4));
			MULT_8_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_8(2,4));
			MULT_8_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_8(2,4));
			MULT_8_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_8(2,4));
			MULT_8_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_8(2,4));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_9(2,4));
			MULT_9_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_9(2,4));
			MULT_9_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_9(2,4));
			MULT_9_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_9(2,4));
			MULT_9_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_9(2,4));
			MULT_9_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_9(2,4));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_10(2,4));
			MULT_10_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_10(2,4));
			MULT_10_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_10(2,4));
			MULT_10_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_10(2,4));
			MULT_10_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_10(2,4));
			MULT_10_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_10(2,4));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_11(2,4));
			MULT_11_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_11(2,4));
			MULT_11_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_11(2,4));
			MULT_11_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_11(2,4));
			MULT_11_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_11(2,4));
			MULT_11_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_11(2,4));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_12(2,4));
			MULT_12_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_12(2,4));
			MULT_12_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_12(2,4));
			MULT_12_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_12(2,4));
			MULT_12_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_12(2,4));
			MULT_12_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_12(2,4));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_13(2,4));
			MULT_13_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_13(2,4));
			MULT_13_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_13(2,4));
			MULT_13_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_13(2,4));
			MULT_13_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_13(2,4));
			MULT_13_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_13(2,4));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_14(2,4));
			MULT_14_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_14(2,4));
			MULT_14_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_14(2,4));
			MULT_14_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_14(2,4));
			MULT_14_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_14(2,4));
			MULT_14_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_14(2,4));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_15(2,4));
			MULT_15_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_15(2,4));
			MULT_15_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_15(2,4));
			MULT_15_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_15(2,4));
			MULT_15_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_15(2,4));
			MULT_15_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_15(2,4));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(2,4)<=signed(WINDOW_1(2,0))*signed(FMAP_1_16(2,4));
			MULT_16_2(2,4)<=signed(WINDOW_2(2,0))*signed(FMAP_2_16(2,4));
			MULT_16_3(2,4)<=signed(WINDOW_3(2,0))*signed(FMAP_3_16(2,4));
			MULT_16_4(2,4)<=signed(WINDOW_4(2,0))*signed(FMAP_4_16(2,4));
			MULT_16_5(2,4)<=signed(WINDOW_5(2,0))*signed(FMAP_5_16(2,4));
			MULT_16_6(2,4)<=signed(WINDOW_6(2,0))*signed(FMAP_6_16(2,4));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(2,4) -----------------------

			MULT_1_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_1(3,0));
			MULT_1_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_1(3,0));
			MULT_1_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_1(3,0));
			MULT_1_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_1(3,0));
			MULT_1_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_1(3,0));
			MULT_1_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_1(3,0));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_2(3,0));
			MULT_2_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_2(3,0));
			MULT_2_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_2(3,0));
			MULT_2_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_2(3,0));
			MULT_2_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_2(3,0));
			MULT_2_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_2(3,0));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_3(3,0));
			MULT_3_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_3(3,0));
			MULT_3_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_3(3,0));
			MULT_3_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_3(3,0));
			MULT_3_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_3(3,0));
			MULT_3_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_3(3,0));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_4(3,0));
			MULT_4_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_4(3,0));
			MULT_4_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_4(3,0));
			MULT_4_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_4(3,0));
			MULT_4_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_4(3,0));
			MULT_4_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_4(3,0));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_5(3,0));
			MULT_5_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_5(3,0));
			MULT_5_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_5(3,0));
			MULT_5_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_5(3,0));
			MULT_5_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_5(3,0));
			MULT_5_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_5(3,0));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_6(3,0));
			MULT_6_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_6(3,0));
			MULT_6_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_6(3,0));
			MULT_6_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_6(3,0));
			MULT_6_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_6(3,0));
			MULT_6_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_6(3,0));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_7(3,0));
			MULT_7_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_7(3,0));
			MULT_7_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_7(3,0));
			MULT_7_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_7(3,0));
			MULT_7_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_7(3,0));
			MULT_7_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_7(3,0));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_8(3,0));
			MULT_8_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_8(3,0));
			MULT_8_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_8(3,0));
			MULT_8_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_8(3,0));
			MULT_8_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_8(3,0));
			MULT_8_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_8(3,0));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_9(3,0));
			MULT_9_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_9(3,0));
			MULT_9_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_9(3,0));
			MULT_9_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_9(3,0));
			MULT_9_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_9(3,0));
			MULT_9_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_9(3,0));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_10(3,0));
			MULT_10_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_10(3,0));
			MULT_10_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_10(3,0));
			MULT_10_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_10(3,0));
			MULT_10_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_10(3,0));
			MULT_10_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_10(3,0));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_11(3,0));
			MULT_11_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_11(3,0));
			MULT_11_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_11(3,0));
			MULT_11_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_11(3,0));
			MULT_11_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_11(3,0));
			MULT_11_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_11(3,0));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_12(3,0));
			MULT_12_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_12(3,0));
			MULT_12_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_12(3,0));
			MULT_12_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_12(3,0));
			MULT_12_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_12(3,0));
			MULT_12_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_12(3,0));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_13(3,0));
			MULT_13_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_13(3,0));
			MULT_13_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_13(3,0));
			MULT_13_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_13(3,0));
			MULT_13_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_13(3,0));
			MULT_13_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_13(3,0));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_14(3,0));
			MULT_14_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_14(3,0));
			MULT_14_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_14(3,0));
			MULT_14_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_14(3,0));
			MULT_14_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_14(3,0));
			MULT_14_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_14(3,0));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_15(3,0));
			MULT_15_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_15(3,0));
			MULT_15_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_15(3,0));
			MULT_15_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_15(3,0));
			MULT_15_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_15(3,0));
			MULT_15_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_15(3,0));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(3,0)<=signed(WINDOW_1(1,4))*signed(FMAP_1_16(3,0));
			MULT_16_2(3,0)<=signed(WINDOW_2(1,4))*signed(FMAP_2_16(3,0));
			MULT_16_3(3,0)<=signed(WINDOW_3(1,4))*signed(FMAP_3_16(3,0));
			MULT_16_4(3,0)<=signed(WINDOW_4(1,4))*signed(FMAP_4_16(3,0));
			MULT_16_5(3,0)<=signed(WINDOW_5(1,4))*signed(FMAP_5_16(3,0));
			MULT_16_6(3,0)<=signed(WINDOW_6(1,4))*signed(FMAP_6_16(3,0));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(3,0) -----------------------

			MULT_1_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_1(3,1));
			MULT_1_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_1(3,1));
			MULT_1_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_1(3,1));
			MULT_1_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_1(3,1));
			MULT_1_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_1(3,1));
			MULT_1_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_1(3,1));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_2(3,1));
			MULT_2_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_2(3,1));
			MULT_2_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_2(3,1));
			MULT_2_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_2(3,1));
			MULT_2_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_2(3,1));
			MULT_2_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_2(3,1));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_3(3,1));
			MULT_3_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_3(3,1));
			MULT_3_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_3(3,1));
			MULT_3_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_3(3,1));
			MULT_3_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_3(3,1));
			MULT_3_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_3(3,1));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_4(3,1));
			MULT_4_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_4(3,1));
			MULT_4_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_4(3,1));
			MULT_4_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_4(3,1));
			MULT_4_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_4(3,1));
			MULT_4_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_4(3,1));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_5(3,1));
			MULT_5_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_5(3,1));
			MULT_5_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_5(3,1));
			MULT_5_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_5(3,1));
			MULT_5_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_5(3,1));
			MULT_5_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_5(3,1));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_6(3,1));
			MULT_6_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_6(3,1));
			MULT_6_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_6(3,1));
			MULT_6_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_6(3,1));
			MULT_6_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_6(3,1));
			MULT_6_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_6(3,1));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_7(3,1));
			MULT_7_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_7(3,1));
			MULT_7_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_7(3,1));
			MULT_7_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_7(3,1));
			MULT_7_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_7(3,1));
			MULT_7_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_7(3,1));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_8(3,1));
			MULT_8_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_8(3,1));
			MULT_8_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_8(3,1));
			MULT_8_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_8(3,1));
			MULT_8_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_8(3,1));
			MULT_8_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_8(3,1));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_9(3,1));
			MULT_9_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_9(3,1));
			MULT_9_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_9(3,1));
			MULT_9_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_9(3,1));
			MULT_9_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_9(3,1));
			MULT_9_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_9(3,1));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_10(3,1));
			MULT_10_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_10(3,1));
			MULT_10_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_10(3,1));
			MULT_10_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_10(3,1));
			MULT_10_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_10(3,1));
			MULT_10_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_10(3,1));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_11(3,1));
			MULT_11_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_11(3,1));
			MULT_11_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_11(3,1));
			MULT_11_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_11(3,1));
			MULT_11_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_11(3,1));
			MULT_11_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_11(3,1));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_12(3,1));
			MULT_12_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_12(3,1));
			MULT_12_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_12(3,1));
			MULT_12_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_12(3,1));
			MULT_12_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_12(3,1));
			MULT_12_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_12(3,1));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_13(3,1));
			MULT_13_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_13(3,1));
			MULT_13_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_13(3,1));
			MULT_13_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_13(3,1));
			MULT_13_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_13(3,1));
			MULT_13_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_13(3,1));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_14(3,1));
			MULT_14_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_14(3,1));
			MULT_14_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_14(3,1));
			MULT_14_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_14(3,1));
			MULT_14_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_14(3,1));
			MULT_14_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_14(3,1));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_15(3,1));
			MULT_15_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_15(3,1));
			MULT_15_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_15(3,1));
			MULT_15_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_15(3,1));
			MULT_15_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_15(3,1));
			MULT_15_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_15(3,1));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(3,1)<=signed(WINDOW_1(1,3))*signed(FMAP_1_16(3,1));
			MULT_16_2(3,1)<=signed(WINDOW_2(1,3))*signed(FMAP_2_16(3,1));
			MULT_16_3(3,1)<=signed(WINDOW_3(1,3))*signed(FMAP_3_16(3,1));
			MULT_16_4(3,1)<=signed(WINDOW_4(1,3))*signed(FMAP_4_16(3,1));
			MULT_16_5(3,1)<=signed(WINDOW_5(1,3))*signed(FMAP_5_16(3,1));
			MULT_16_6(3,1)<=signed(WINDOW_6(1,3))*signed(FMAP_6_16(3,1));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(3,1) -----------------------

			MULT_1_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_1(3,2));
			MULT_1_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_1(3,2));
			MULT_1_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_1(3,2));
			MULT_1_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_1(3,2));
			MULT_1_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_1(3,2));
			MULT_1_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_1(3,2));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_2(3,2));
			MULT_2_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_2(3,2));
			MULT_2_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_2(3,2));
			MULT_2_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_2(3,2));
			MULT_2_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_2(3,2));
			MULT_2_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_2(3,2));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_3(3,2));
			MULT_3_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_3(3,2));
			MULT_3_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_3(3,2));
			MULT_3_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_3(3,2));
			MULT_3_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_3(3,2));
			MULT_3_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_3(3,2));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_4(3,2));
			MULT_4_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_4(3,2));
			MULT_4_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_4(3,2));
			MULT_4_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_4(3,2));
			MULT_4_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_4(3,2));
			MULT_4_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_4(3,2));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_5(3,2));
			MULT_5_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_5(3,2));
			MULT_5_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_5(3,2));
			MULT_5_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_5(3,2));
			MULT_5_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_5(3,2));
			MULT_5_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_5(3,2));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_6(3,2));
			MULT_6_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_6(3,2));
			MULT_6_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_6(3,2));
			MULT_6_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_6(3,2));
			MULT_6_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_6(3,2));
			MULT_6_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_6(3,2));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_7(3,2));
			MULT_7_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_7(3,2));
			MULT_7_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_7(3,2));
			MULT_7_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_7(3,2));
			MULT_7_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_7(3,2));
			MULT_7_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_7(3,2));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_8(3,2));
			MULT_8_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_8(3,2));
			MULT_8_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_8(3,2));
			MULT_8_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_8(3,2));
			MULT_8_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_8(3,2));
			MULT_8_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_8(3,2));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_9(3,2));
			MULT_9_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_9(3,2));
			MULT_9_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_9(3,2));
			MULT_9_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_9(3,2));
			MULT_9_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_9(3,2));
			MULT_9_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_9(3,2));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_10(3,2));
			MULT_10_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_10(3,2));
			MULT_10_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_10(3,2));
			MULT_10_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_10(3,2));
			MULT_10_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_10(3,2));
			MULT_10_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_10(3,2));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_11(3,2));
			MULT_11_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_11(3,2));
			MULT_11_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_11(3,2));
			MULT_11_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_11(3,2));
			MULT_11_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_11(3,2));
			MULT_11_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_11(3,2));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_12(3,2));
			MULT_12_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_12(3,2));
			MULT_12_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_12(3,2));
			MULT_12_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_12(3,2));
			MULT_12_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_12(3,2));
			MULT_12_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_12(3,2));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_13(3,2));
			MULT_13_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_13(3,2));
			MULT_13_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_13(3,2));
			MULT_13_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_13(3,2));
			MULT_13_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_13(3,2));
			MULT_13_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_13(3,2));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_14(3,2));
			MULT_14_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_14(3,2));
			MULT_14_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_14(3,2));
			MULT_14_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_14(3,2));
			MULT_14_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_14(3,2));
			MULT_14_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_14(3,2));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_15(3,2));
			MULT_15_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_15(3,2));
			MULT_15_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_15(3,2));
			MULT_15_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_15(3,2));
			MULT_15_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_15(3,2));
			MULT_15_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_15(3,2));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(3,2)<=signed(WINDOW_1(1,2))*signed(FMAP_1_16(3,2));
			MULT_16_2(3,2)<=signed(WINDOW_2(1,2))*signed(FMAP_2_16(3,2));
			MULT_16_3(3,2)<=signed(WINDOW_3(1,2))*signed(FMAP_3_16(3,2));
			MULT_16_4(3,2)<=signed(WINDOW_4(1,2))*signed(FMAP_4_16(3,2));
			MULT_16_5(3,2)<=signed(WINDOW_5(1,2))*signed(FMAP_5_16(3,2));
			MULT_16_6(3,2)<=signed(WINDOW_6(1,2))*signed(FMAP_6_16(3,2));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(3,2) -----------------------

			MULT_1_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_1(3,3));
			MULT_1_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_1(3,3));
			MULT_1_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_1(3,3));
			MULT_1_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_1(3,3));
			MULT_1_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_1(3,3));
			MULT_1_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_1(3,3));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_2(3,3));
			MULT_2_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_2(3,3));
			MULT_2_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_2(3,3));
			MULT_2_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_2(3,3));
			MULT_2_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_2(3,3));
			MULT_2_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_2(3,3));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_3(3,3));
			MULT_3_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_3(3,3));
			MULT_3_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_3(3,3));
			MULT_3_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_3(3,3));
			MULT_3_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_3(3,3));
			MULT_3_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_3(3,3));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_4(3,3));
			MULT_4_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_4(3,3));
			MULT_4_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_4(3,3));
			MULT_4_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_4(3,3));
			MULT_4_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_4(3,3));
			MULT_4_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_4(3,3));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_5(3,3));
			MULT_5_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_5(3,3));
			MULT_5_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_5(3,3));
			MULT_5_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_5(3,3));
			MULT_5_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_5(3,3));
			MULT_5_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_5(3,3));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_6(3,3));
			MULT_6_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_6(3,3));
			MULT_6_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_6(3,3));
			MULT_6_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_6(3,3));
			MULT_6_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_6(3,3));
			MULT_6_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_6(3,3));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_7(3,3));
			MULT_7_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_7(3,3));
			MULT_7_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_7(3,3));
			MULT_7_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_7(3,3));
			MULT_7_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_7(3,3));
			MULT_7_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_7(3,3));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_8(3,3));
			MULT_8_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_8(3,3));
			MULT_8_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_8(3,3));
			MULT_8_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_8(3,3));
			MULT_8_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_8(3,3));
			MULT_8_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_8(3,3));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_9(3,3));
			MULT_9_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_9(3,3));
			MULT_9_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_9(3,3));
			MULT_9_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_9(3,3));
			MULT_9_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_9(3,3));
			MULT_9_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_9(3,3));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_10(3,3));
			MULT_10_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_10(3,3));
			MULT_10_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_10(3,3));
			MULT_10_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_10(3,3));
			MULT_10_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_10(3,3));
			MULT_10_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_10(3,3));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_11(3,3));
			MULT_11_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_11(3,3));
			MULT_11_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_11(3,3));
			MULT_11_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_11(3,3));
			MULT_11_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_11(3,3));
			MULT_11_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_11(3,3));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_12(3,3));
			MULT_12_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_12(3,3));
			MULT_12_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_12(3,3));
			MULT_12_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_12(3,3));
			MULT_12_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_12(3,3));
			MULT_12_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_12(3,3));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_13(3,3));
			MULT_13_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_13(3,3));
			MULT_13_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_13(3,3));
			MULT_13_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_13(3,3));
			MULT_13_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_13(3,3));
			MULT_13_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_13(3,3));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_14(3,3));
			MULT_14_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_14(3,3));
			MULT_14_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_14(3,3));
			MULT_14_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_14(3,3));
			MULT_14_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_14(3,3));
			MULT_14_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_14(3,3));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_15(3,3));
			MULT_15_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_15(3,3));
			MULT_15_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_15(3,3));
			MULT_15_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_15(3,3));
			MULT_15_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_15(3,3));
			MULT_15_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_15(3,3));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(3,3)<=signed(WINDOW_1(1,1))*signed(FMAP_1_16(3,3));
			MULT_16_2(3,3)<=signed(WINDOW_2(1,1))*signed(FMAP_2_16(3,3));
			MULT_16_3(3,3)<=signed(WINDOW_3(1,1))*signed(FMAP_3_16(3,3));
			MULT_16_4(3,3)<=signed(WINDOW_4(1,1))*signed(FMAP_4_16(3,3));
			MULT_16_5(3,3)<=signed(WINDOW_5(1,1))*signed(FMAP_5_16(3,3));
			MULT_16_6(3,3)<=signed(WINDOW_6(1,1))*signed(FMAP_6_16(3,3));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(3,3) -----------------------

			MULT_1_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_1(3,4));
			MULT_1_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_1(3,4));
			MULT_1_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_1(3,4));
			MULT_1_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_1(3,4));
			MULT_1_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_1(3,4));
			MULT_1_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_1(3,4));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_2(3,4));
			MULT_2_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_2(3,4));
			MULT_2_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_2(3,4));
			MULT_2_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_2(3,4));
			MULT_2_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_2(3,4));
			MULT_2_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_2(3,4));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_3(3,4));
			MULT_3_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_3(3,4));
			MULT_3_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_3(3,4));
			MULT_3_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_3(3,4));
			MULT_3_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_3(3,4));
			MULT_3_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_3(3,4));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_4(3,4));
			MULT_4_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_4(3,4));
			MULT_4_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_4(3,4));
			MULT_4_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_4(3,4));
			MULT_4_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_4(3,4));
			MULT_4_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_4(3,4));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_5(3,4));
			MULT_5_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_5(3,4));
			MULT_5_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_5(3,4));
			MULT_5_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_5(3,4));
			MULT_5_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_5(3,4));
			MULT_5_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_5(3,4));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_6(3,4));
			MULT_6_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_6(3,4));
			MULT_6_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_6(3,4));
			MULT_6_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_6(3,4));
			MULT_6_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_6(3,4));
			MULT_6_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_6(3,4));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_7(3,4));
			MULT_7_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_7(3,4));
			MULT_7_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_7(3,4));
			MULT_7_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_7(3,4));
			MULT_7_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_7(3,4));
			MULT_7_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_7(3,4));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_8(3,4));
			MULT_8_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_8(3,4));
			MULT_8_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_8(3,4));
			MULT_8_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_8(3,4));
			MULT_8_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_8(3,4));
			MULT_8_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_8(3,4));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_9(3,4));
			MULT_9_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_9(3,4));
			MULT_9_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_9(3,4));
			MULT_9_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_9(3,4));
			MULT_9_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_9(3,4));
			MULT_9_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_9(3,4));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_10(3,4));
			MULT_10_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_10(3,4));
			MULT_10_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_10(3,4));
			MULT_10_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_10(3,4));
			MULT_10_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_10(3,4));
			MULT_10_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_10(3,4));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_11(3,4));
			MULT_11_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_11(3,4));
			MULT_11_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_11(3,4));
			MULT_11_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_11(3,4));
			MULT_11_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_11(3,4));
			MULT_11_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_11(3,4));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_12(3,4));
			MULT_12_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_12(3,4));
			MULT_12_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_12(3,4));
			MULT_12_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_12(3,4));
			MULT_12_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_12(3,4));
			MULT_12_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_12(3,4));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_13(3,4));
			MULT_13_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_13(3,4));
			MULT_13_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_13(3,4));
			MULT_13_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_13(3,4));
			MULT_13_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_13(3,4));
			MULT_13_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_13(3,4));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_14(3,4));
			MULT_14_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_14(3,4));
			MULT_14_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_14(3,4));
			MULT_14_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_14(3,4));
			MULT_14_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_14(3,4));
			MULT_14_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_14(3,4));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_15(3,4));
			MULT_15_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_15(3,4));
			MULT_15_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_15(3,4));
			MULT_15_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_15(3,4));
			MULT_15_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_15(3,4));
			MULT_15_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_15(3,4));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(3,4)<=signed(WINDOW_1(1,0))*signed(FMAP_1_16(3,4));
			MULT_16_2(3,4)<=signed(WINDOW_2(1,0))*signed(FMAP_2_16(3,4));
			MULT_16_3(3,4)<=signed(WINDOW_3(1,0))*signed(FMAP_3_16(3,4));
			MULT_16_4(3,4)<=signed(WINDOW_4(1,0))*signed(FMAP_4_16(3,4));
			MULT_16_5(3,4)<=signed(WINDOW_5(1,0))*signed(FMAP_5_16(3,4));
			MULT_16_6(3,4)<=signed(WINDOW_6(1,0))*signed(FMAP_6_16(3,4));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(3,4) -----------------------

			MULT_1_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_1(4,0));
			MULT_1_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_1(4,0));
			MULT_1_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_1(4,0));
			MULT_1_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_1(4,0));
			MULT_1_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_1(4,0));
			MULT_1_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_1(4,0));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_2(4,0));
			MULT_2_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_2(4,0));
			MULT_2_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_2(4,0));
			MULT_2_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_2(4,0));
			MULT_2_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_2(4,0));
			MULT_2_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_2(4,0));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_3(4,0));
			MULT_3_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_3(4,0));
			MULT_3_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_3(4,0));
			MULT_3_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_3(4,0));
			MULT_3_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_3(4,0));
			MULT_3_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_3(4,0));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_4(4,0));
			MULT_4_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_4(4,0));
			MULT_4_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_4(4,0));
			MULT_4_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_4(4,0));
			MULT_4_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_4(4,0));
			MULT_4_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_4(4,0));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_5(4,0));
			MULT_5_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_5(4,0));
			MULT_5_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_5(4,0));
			MULT_5_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_5(4,0));
			MULT_5_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_5(4,0));
			MULT_5_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_5(4,0));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_6(4,0));
			MULT_6_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_6(4,0));
			MULT_6_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_6(4,0));
			MULT_6_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_6(4,0));
			MULT_6_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_6(4,0));
			MULT_6_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_6(4,0));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_7(4,0));
			MULT_7_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_7(4,0));
			MULT_7_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_7(4,0));
			MULT_7_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_7(4,0));
			MULT_7_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_7(4,0));
			MULT_7_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_7(4,0));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_8(4,0));
			MULT_8_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_8(4,0));
			MULT_8_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_8(4,0));
			MULT_8_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_8(4,0));
			MULT_8_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_8(4,0));
			MULT_8_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_8(4,0));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_9(4,0));
			MULT_9_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_9(4,0));
			MULT_9_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_9(4,0));
			MULT_9_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_9(4,0));
			MULT_9_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_9(4,0));
			MULT_9_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_9(4,0));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_10(4,0));
			MULT_10_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_10(4,0));
			MULT_10_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_10(4,0));
			MULT_10_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_10(4,0));
			MULT_10_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_10(4,0));
			MULT_10_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_10(4,0));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_11(4,0));
			MULT_11_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_11(4,0));
			MULT_11_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_11(4,0));
			MULT_11_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_11(4,0));
			MULT_11_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_11(4,0));
			MULT_11_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_11(4,0));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_12(4,0));
			MULT_12_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_12(4,0));
			MULT_12_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_12(4,0));
			MULT_12_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_12(4,0));
			MULT_12_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_12(4,0));
			MULT_12_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_12(4,0));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_13(4,0));
			MULT_13_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_13(4,0));
			MULT_13_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_13(4,0));
			MULT_13_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_13(4,0));
			MULT_13_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_13(4,0));
			MULT_13_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_13(4,0));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_14(4,0));
			MULT_14_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_14(4,0));
			MULT_14_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_14(4,0));
			MULT_14_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_14(4,0));
			MULT_14_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_14(4,0));
			MULT_14_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_14(4,0));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_15(4,0));
			MULT_15_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_15(4,0));
			MULT_15_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_15(4,0));
			MULT_15_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_15(4,0));
			MULT_15_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_15(4,0));
			MULT_15_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_15(4,0));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(4,0)<=signed(WINDOW_1(0,4))*signed(FMAP_1_16(4,0));
			MULT_16_2(4,0)<=signed(WINDOW_2(0,4))*signed(FMAP_2_16(4,0));
			MULT_16_3(4,0)<=signed(WINDOW_3(0,4))*signed(FMAP_3_16(4,0));
			MULT_16_4(4,0)<=signed(WINDOW_4(0,4))*signed(FMAP_4_16(4,0));
			MULT_16_5(4,0)<=signed(WINDOW_5(0,4))*signed(FMAP_5_16(4,0));
			MULT_16_6(4,0)<=signed(WINDOW_6(0,4))*signed(FMAP_6_16(4,0));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(4,0) -----------------------

			MULT_1_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_1(4,1));
			MULT_1_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_1(4,1));
			MULT_1_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_1(4,1));
			MULT_1_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_1(4,1));
			MULT_1_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_1(4,1));
			MULT_1_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_1(4,1));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_2(4,1));
			MULT_2_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_2(4,1));
			MULT_2_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_2(4,1));
			MULT_2_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_2(4,1));
			MULT_2_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_2(4,1));
			MULT_2_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_2(4,1));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_3(4,1));
			MULT_3_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_3(4,1));
			MULT_3_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_3(4,1));
			MULT_3_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_3(4,1));
			MULT_3_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_3(4,1));
			MULT_3_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_3(4,1));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_4(4,1));
			MULT_4_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_4(4,1));
			MULT_4_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_4(4,1));
			MULT_4_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_4(4,1));
			MULT_4_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_4(4,1));
			MULT_4_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_4(4,1));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_5(4,1));
			MULT_5_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_5(4,1));
			MULT_5_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_5(4,1));
			MULT_5_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_5(4,1));
			MULT_5_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_5(4,1));
			MULT_5_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_5(4,1));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_6(4,1));
			MULT_6_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_6(4,1));
			MULT_6_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_6(4,1));
			MULT_6_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_6(4,1));
			MULT_6_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_6(4,1));
			MULT_6_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_6(4,1));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_7(4,1));
			MULT_7_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_7(4,1));
			MULT_7_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_7(4,1));
			MULT_7_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_7(4,1));
			MULT_7_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_7(4,1));
			MULT_7_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_7(4,1));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_8(4,1));
			MULT_8_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_8(4,1));
			MULT_8_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_8(4,1));
			MULT_8_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_8(4,1));
			MULT_8_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_8(4,1));
			MULT_8_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_8(4,1));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_9(4,1));
			MULT_9_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_9(4,1));
			MULT_9_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_9(4,1));
			MULT_9_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_9(4,1));
			MULT_9_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_9(4,1));
			MULT_9_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_9(4,1));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_10(4,1));
			MULT_10_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_10(4,1));
			MULT_10_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_10(4,1));
			MULT_10_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_10(4,1));
			MULT_10_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_10(4,1));
			MULT_10_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_10(4,1));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_11(4,1));
			MULT_11_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_11(4,1));
			MULT_11_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_11(4,1));
			MULT_11_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_11(4,1));
			MULT_11_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_11(4,1));
			MULT_11_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_11(4,1));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_12(4,1));
			MULT_12_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_12(4,1));
			MULT_12_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_12(4,1));
			MULT_12_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_12(4,1));
			MULT_12_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_12(4,1));
			MULT_12_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_12(4,1));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_13(4,1));
			MULT_13_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_13(4,1));
			MULT_13_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_13(4,1));
			MULT_13_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_13(4,1));
			MULT_13_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_13(4,1));
			MULT_13_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_13(4,1));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_14(4,1));
			MULT_14_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_14(4,1));
			MULT_14_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_14(4,1));
			MULT_14_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_14(4,1));
			MULT_14_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_14(4,1));
			MULT_14_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_14(4,1));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_15(4,1));
			MULT_15_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_15(4,1));
			MULT_15_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_15(4,1));
			MULT_15_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_15(4,1));
			MULT_15_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_15(4,1));
			MULT_15_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_15(4,1));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(4,1)<=signed(WINDOW_1(0,3))*signed(FMAP_1_16(4,1));
			MULT_16_2(4,1)<=signed(WINDOW_2(0,3))*signed(FMAP_2_16(4,1));
			MULT_16_3(4,1)<=signed(WINDOW_3(0,3))*signed(FMAP_3_16(4,1));
			MULT_16_4(4,1)<=signed(WINDOW_4(0,3))*signed(FMAP_4_16(4,1));
			MULT_16_5(4,1)<=signed(WINDOW_5(0,3))*signed(FMAP_5_16(4,1));
			MULT_16_6(4,1)<=signed(WINDOW_6(0,3))*signed(FMAP_6_16(4,1));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(4,1) -----------------------

			MULT_1_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_1(4,2));
			MULT_1_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_1(4,2));
			MULT_1_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_1(4,2));
			MULT_1_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_1(4,2));
			MULT_1_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_1(4,2));
			MULT_1_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_1(4,2));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_2(4,2));
			MULT_2_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_2(4,2));
			MULT_2_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_2(4,2));
			MULT_2_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_2(4,2));
			MULT_2_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_2(4,2));
			MULT_2_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_2(4,2));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_3(4,2));
			MULT_3_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_3(4,2));
			MULT_3_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_3(4,2));
			MULT_3_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_3(4,2));
			MULT_3_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_3(4,2));
			MULT_3_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_3(4,2));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_4(4,2));
			MULT_4_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_4(4,2));
			MULT_4_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_4(4,2));
			MULT_4_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_4(4,2));
			MULT_4_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_4(4,2));
			MULT_4_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_4(4,2));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_5(4,2));
			MULT_5_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_5(4,2));
			MULT_5_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_5(4,2));
			MULT_5_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_5(4,2));
			MULT_5_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_5(4,2));
			MULT_5_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_5(4,2));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_6(4,2));
			MULT_6_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_6(4,2));
			MULT_6_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_6(4,2));
			MULT_6_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_6(4,2));
			MULT_6_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_6(4,2));
			MULT_6_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_6(4,2));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_7(4,2));
			MULT_7_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_7(4,2));
			MULT_7_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_7(4,2));
			MULT_7_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_7(4,2));
			MULT_7_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_7(4,2));
			MULT_7_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_7(4,2));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_8(4,2));
			MULT_8_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_8(4,2));
			MULT_8_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_8(4,2));
			MULT_8_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_8(4,2));
			MULT_8_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_8(4,2));
			MULT_8_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_8(4,2));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_9(4,2));
			MULT_9_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_9(4,2));
			MULT_9_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_9(4,2));
			MULT_9_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_9(4,2));
			MULT_9_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_9(4,2));
			MULT_9_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_9(4,2));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_10(4,2));
			MULT_10_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_10(4,2));
			MULT_10_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_10(4,2));
			MULT_10_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_10(4,2));
			MULT_10_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_10(4,2));
			MULT_10_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_10(4,2));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_11(4,2));
			MULT_11_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_11(4,2));
			MULT_11_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_11(4,2));
			MULT_11_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_11(4,2));
			MULT_11_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_11(4,2));
			MULT_11_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_11(4,2));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_12(4,2));
			MULT_12_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_12(4,2));
			MULT_12_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_12(4,2));
			MULT_12_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_12(4,2));
			MULT_12_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_12(4,2));
			MULT_12_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_12(4,2));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_13(4,2));
			MULT_13_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_13(4,2));
			MULT_13_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_13(4,2));
			MULT_13_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_13(4,2));
			MULT_13_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_13(4,2));
			MULT_13_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_13(4,2));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_14(4,2));
			MULT_14_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_14(4,2));
			MULT_14_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_14(4,2));
			MULT_14_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_14(4,2));
			MULT_14_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_14(4,2));
			MULT_14_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_14(4,2));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_15(4,2));
			MULT_15_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_15(4,2));
			MULT_15_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_15(4,2));
			MULT_15_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_15(4,2));
			MULT_15_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_15(4,2));
			MULT_15_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_15(4,2));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(4,2)<=signed(WINDOW_1(0,2))*signed(FMAP_1_16(4,2));
			MULT_16_2(4,2)<=signed(WINDOW_2(0,2))*signed(FMAP_2_16(4,2));
			MULT_16_3(4,2)<=signed(WINDOW_3(0,2))*signed(FMAP_3_16(4,2));
			MULT_16_4(4,2)<=signed(WINDOW_4(0,2))*signed(FMAP_4_16(4,2));
			MULT_16_5(4,2)<=signed(WINDOW_5(0,2))*signed(FMAP_5_16(4,2));
			MULT_16_6(4,2)<=signed(WINDOW_6(0,2))*signed(FMAP_6_16(4,2));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(4,2) -----------------------

			MULT_1_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_1(4,3));
			MULT_1_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_1(4,3));
			MULT_1_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_1(4,3));
			MULT_1_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_1(4,3));
			MULT_1_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_1(4,3));
			MULT_1_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_1(4,3));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_2(4,3));
			MULT_2_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_2(4,3));
			MULT_2_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_2(4,3));
			MULT_2_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_2(4,3));
			MULT_2_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_2(4,3));
			MULT_2_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_2(4,3));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_3(4,3));
			MULT_3_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_3(4,3));
			MULT_3_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_3(4,3));
			MULT_3_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_3(4,3));
			MULT_3_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_3(4,3));
			MULT_3_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_3(4,3));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_4(4,3));
			MULT_4_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_4(4,3));
			MULT_4_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_4(4,3));
			MULT_4_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_4(4,3));
			MULT_4_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_4(4,3));
			MULT_4_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_4(4,3));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_5(4,3));
			MULT_5_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_5(4,3));
			MULT_5_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_5(4,3));
			MULT_5_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_5(4,3));
			MULT_5_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_5(4,3));
			MULT_5_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_5(4,3));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_6(4,3));
			MULT_6_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_6(4,3));
			MULT_6_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_6(4,3));
			MULT_6_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_6(4,3));
			MULT_6_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_6(4,3));
			MULT_6_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_6(4,3));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_7(4,3));
			MULT_7_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_7(4,3));
			MULT_7_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_7(4,3));
			MULT_7_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_7(4,3));
			MULT_7_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_7(4,3));
			MULT_7_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_7(4,3));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_8(4,3));
			MULT_8_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_8(4,3));
			MULT_8_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_8(4,3));
			MULT_8_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_8(4,3));
			MULT_8_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_8(4,3));
			MULT_8_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_8(4,3));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_9(4,3));
			MULT_9_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_9(4,3));
			MULT_9_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_9(4,3));
			MULT_9_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_9(4,3));
			MULT_9_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_9(4,3));
			MULT_9_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_9(4,3));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_10(4,3));
			MULT_10_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_10(4,3));
			MULT_10_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_10(4,3));
			MULT_10_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_10(4,3));
			MULT_10_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_10(4,3));
			MULT_10_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_10(4,3));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_11(4,3));
			MULT_11_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_11(4,3));
			MULT_11_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_11(4,3));
			MULT_11_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_11(4,3));
			MULT_11_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_11(4,3));
			MULT_11_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_11(4,3));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_12(4,3));
			MULT_12_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_12(4,3));
			MULT_12_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_12(4,3));
			MULT_12_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_12(4,3));
			MULT_12_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_12(4,3));
			MULT_12_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_12(4,3));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_13(4,3));
			MULT_13_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_13(4,3));
			MULT_13_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_13(4,3));
			MULT_13_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_13(4,3));
			MULT_13_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_13(4,3));
			MULT_13_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_13(4,3));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_14(4,3));
			MULT_14_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_14(4,3));
			MULT_14_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_14(4,3));
			MULT_14_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_14(4,3));
			MULT_14_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_14(4,3));
			MULT_14_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_14(4,3));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_15(4,3));
			MULT_15_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_15(4,3));
			MULT_15_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_15(4,3));
			MULT_15_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_15(4,3));
			MULT_15_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_15(4,3));
			MULT_15_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_15(4,3));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(4,3)<=signed(WINDOW_1(0,1))*signed(FMAP_1_16(4,3));
			MULT_16_2(4,3)<=signed(WINDOW_2(0,1))*signed(FMAP_2_16(4,3));
			MULT_16_3(4,3)<=signed(WINDOW_3(0,1))*signed(FMAP_3_16(4,3));
			MULT_16_4(4,3)<=signed(WINDOW_4(0,1))*signed(FMAP_4_16(4,3));
			MULT_16_5(4,3)<=signed(WINDOW_5(0,1))*signed(FMAP_5_16(4,3));
			MULT_16_6(4,3)<=signed(WINDOW_6(0,1))*signed(FMAP_6_16(4,3));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(4,3) -----------------------

			MULT_1_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_1(4,4));
			MULT_1_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_1(4,4));
			MULT_1_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_1(4,4));
			MULT_1_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_1(4,4));
			MULT_1_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_1(4,4));
			MULT_1_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_1(4,4));
			------------------------- END FMAP(1) ---------------------
			MULT_2_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_2(4,4));
			MULT_2_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_2(4,4));
			MULT_2_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_2(4,4));
			MULT_2_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_2(4,4));
			MULT_2_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_2(4,4));
			MULT_2_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_2(4,4));
			------------------------- END FMAP(2) ---------------------
			MULT_3_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_3(4,4));
			MULT_3_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_3(4,4));
			MULT_3_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_3(4,4));
			MULT_3_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_3(4,4));
			MULT_3_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_3(4,4));
			MULT_3_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_3(4,4));
			------------------------- END FMAP(3) ---------------------
			MULT_4_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_4(4,4));
			MULT_4_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_4(4,4));
			MULT_4_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_4(4,4));
			MULT_4_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_4(4,4));
			MULT_4_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_4(4,4));
			MULT_4_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_4(4,4));
			------------------------- END FMAP(4) ---------------------
			MULT_5_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_5(4,4));
			MULT_5_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_5(4,4));
			MULT_5_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_5(4,4));
			MULT_5_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_5(4,4));
			MULT_5_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_5(4,4));
			MULT_5_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_5(4,4));
			------------------------- END FMAP(5) ---------------------
			MULT_6_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_6(4,4));
			MULT_6_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_6(4,4));
			MULT_6_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_6(4,4));
			MULT_6_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_6(4,4));
			MULT_6_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_6(4,4));
			MULT_6_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_6(4,4));
			------------------------- END FMAP(6) ---------------------
			MULT_7_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_7(4,4));
			MULT_7_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_7(4,4));
			MULT_7_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_7(4,4));
			MULT_7_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_7(4,4));
			MULT_7_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_7(4,4));
			MULT_7_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_7(4,4));
			------------------------- END FMAP(7) ---------------------
			MULT_8_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_8(4,4));
			MULT_8_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_8(4,4));
			MULT_8_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_8(4,4));
			MULT_8_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_8(4,4));
			MULT_8_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_8(4,4));
			MULT_8_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_8(4,4));
			------------------------- END FMAP(8) ---------------------
			MULT_9_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_9(4,4));
			MULT_9_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_9(4,4));
			MULT_9_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_9(4,4));
			MULT_9_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_9(4,4));
			MULT_9_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_9(4,4));
			MULT_9_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_9(4,4));
			------------------------- END FMAP(9) ---------------------
			MULT_10_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_10(4,4));
			MULT_10_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_10(4,4));
			MULT_10_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_10(4,4));
			MULT_10_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_10(4,4));
			MULT_10_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_10(4,4));
			MULT_10_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_10(4,4));
			------------------------- END FMAP(10) ---------------------
			MULT_11_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_11(4,4));
			MULT_11_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_11(4,4));
			MULT_11_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_11(4,4));
			MULT_11_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_11(4,4));
			MULT_11_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_11(4,4));
			MULT_11_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_11(4,4));
			------------------------- END FMAP(11) ---------------------
			MULT_12_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_12(4,4));
			MULT_12_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_12(4,4));
			MULT_12_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_12(4,4));
			MULT_12_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_12(4,4));
			MULT_12_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_12(4,4));
			MULT_12_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_12(4,4));
			------------------------- END FMAP(12) ---------------------
			MULT_13_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_13(4,4));
			MULT_13_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_13(4,4));
			MULT_13_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_13(4,4));
			MULT_13_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_13(4,4));
			MULT_13_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_13(4,4));
			MULT_13_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_13(4,4));
			------------------------- END FMAP(13) ---------------------
			MULT_14_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_14(4,4));
			MULT_14_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_14(4,4));
			MULT_14_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_14(4,4));
			MULT_14_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_14(4,4));
			MULT_14_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_14(4,4));
			MULT_14_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_14(4,4));
			------------------------- END FMAP(14) ---------------------
			MULT_15_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_15(4,4));
			MULT_15_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_15(4,4));
			MULT_15_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_15(4,4));
			MULT_15_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_15(4,4));
			MULT_15_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_15(4,4));
			MULT_15_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_15(4,4));
			------------------------- END FMAP(15) ---------------------
			MULT_16_1(4,4)<=signed(WINDOW_1(0,0))*signed(FMAP_1_16(4,4));
			MULT_16_2(4,4)<=signed(WINDOW_2(0,0))*signed(FMAP_2_16(4,4));
			MULT_16_3(4,4)<=signed(WINDOW_3(0,0))*signed(FMAP_3_16(4,4));
			MULT_16_4(4,4)<=signed(WINDOW_4(0,0))*signed(FMAP_4_16(4,4));
			MULT_16_5(4,4)<=signed(WINDOW_5(0,0))*signed(FMAP_5_16(4,4));
			MULT_16_6(4,4)<=signed(WINDOW_6(0,0))*signed(FMAP_6_16(4,4));
			------------------------- END FMAP(16) ---------------------
			-------------------------END OF INDEX(4,4) -----------------------


			EN_SUM_MULT_1<='1';	
		end if;

		------------------------- Enable SUM_MULT START -----------------------
		if EN_SUM_MULT_1 = '1' then
			------------------------------------STAGE-1--------------------------------------
			MULTS_1_1_1(0,0)<=signed(MULT_1_1(0,0)(MULT_SIZE-1) & MULT_1_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(0,0)(MULT_SIZE-1) & MULT_1_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(0,0)<=signed(MULT_1_3(0,0)(MULT_SIZE-1) & MULT_1_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(0,0)(MULT_SIZE-1) & MULT_1_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(0,0)<=signed(MULT_1_5(0,0)(MULT_SIZE-1) & MULT_1_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(0,0)(MULT_SIZE-1) & MULT_1_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(0,0)<=signed(MULT_2_1(0,0)(MULT_SIZE-1) & MULT_2_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(0,0)(MULT_SIZE-1) & MULT_2_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(0,0)<=signed(MULT_2_3(0,0)(MULT_SIZE-1) & MULT_2_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(0,0)(MULT_SIZE-1) & MULT_2_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(0,0)<=signed(MULT_2_5(0,0)(MULT_SIZE-1) & MULT_2_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(0,0)(MULT_SIZE-1) & MULT_2_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(0,0)<=signed(MULT_3_1(0,0)(MULT_SIZE-1) & MULT_3_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(0,0)(MULT_SIZE-1) & MULT_3_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(0,0)<=signed(MULT_3_3(0,0)(MULT_SIZE-1) & MULT_3_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(0,0)(MULT_SIZE-1) & MULT_3_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(0,0)<=signed(MULT_3_5(0,0)(MULT_SIZE-1) & MULT_3_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(0,0)(MULT_SIZE-1) & MULT_3_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(0,0)<=signed(MULT_4_1(0,0)(MULT_SIZE-1) & MULT_4_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(0,0)(MULT_SIZE-1) & MULT_4_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(0,0)<=signed(MULT_4_3(0,0)(MULT_SIZE-1) & MULT_4_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(0,0)(MULT_SIZE-1) & MULT_4_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(0,0)<=signed(MULT_4_5(0,0)(MULT_SIZE-1) & MULT_4_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(0,0)(MULT_SIZE-1) & MULT_4_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(0,0)<=signed(MULT_5_1(0,0)(MULT_SIZE-1) & MULT_5_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(0,0)(MULT_SIZE-1) & MULT_5_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(0,0)<=signed(MULT_5_3(0,0)(MULT_SIZE-1) & MULT_5_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(0,0)(MULT_SIZE-1) & MULT_5_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(0,0)<=signed(MULT_5_5(0,0)(MULT_SIZE-1) & MULT_5_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(0,0)(MULT_SIZE-1) & MULT_5_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(0,0)<=signed(MULT_6_1(0,0)(MULT_SIZE-1) & MULT_6_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(0,0)(MULT_SIZE-1) & MULT_6_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(0,0)<=signed(MULT_6_3(0,0)(MULT_SIZE-1) & MULT_6_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(0,0)(MULT_SIZE-1) & MULT_6_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(0,0)<=signed(MULT_6_5(0,0)(MULT_SIZE-1) & MULT_6_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(0,0)(MULT_SIZE-1) & MULT_6_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(0,0)<=signed(MULT_7_1(0,0)(MULT_SIZE-1) & MULT_7_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(0,0)(MULT_SIZE-1) & MULT_7_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(0,0)<=signed(MULT_7_3(0,0)(MULT_SIZE-1) & MULT_7_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(0,0)(MULT_SIZE-1) & MULT_7_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(0,0)<=signed(MULT_7_5(0,0)(MULT_SIZE-1) & MULT_7_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(0,0)(MULT_SIZE-1) & MULT_7_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(0,0)<=signed(MULT_8_1(0,0)(MULT_SIZE-1) & MULT_8_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(0,0)(MULT_SIZE-1) & MULT_8_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(0,0)<=signed(MULT_8_3(0,0)(MULT_SIZE-1) & MULT_8_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(0,0)(MULT_SIZE-1) & MULT_8_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(0,0)<=signed(MULT_8_5(0,0)(MULT_SIZE-1) & MULT_8_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(0,0)(MULT_SIZE-1) & MULT_8_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(0,0)<=signed(MULT_9_1(0,0)(MULT_SIZE-1) & MULT_9_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(0,0)(MULT_SIZE-1) & MULT_9_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(0,0)<=signed(MULT_9_3(0,0)(MULT_SIZE-1) & MULT_9_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(0,0)(MULT_SIZE-1) & MULT_9_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(0,0)<=signed(MULT_9_5(0,0)(MULT_SIZE-1) & MULT_9_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(0,0)(MULT_SIZE-1) & MULT_9_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(0,0)<=signed(MULT_10_1(0,0)(MULT_SIZE-1) & MULT_10_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(0,0)(MULT_SIZE-1) & MULT_10_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(0,0)<=signed(MULT_10_3(0,0)(MULT_SIZE-1) & MULT_10_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(0,0)(MULT_SIZE-1) & MULT_10_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(0,0)<=signed(MULT_10_5(0,0)(MULT_SIZE-1) & MULT_10_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(0,0)(MULT_SIZE-1) & MULT_10_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(0,0)<=signed(MULT_11_1(0,0)(MULT_SIZE-1) & MULT_11_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(0,0)(MULT_SIZE-1) & MULT_11_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(0,0)<=signed(MULT_11_3(0,0)(MULT_SIZE-1) & MULT_11_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(0,0)(MULT_SIZE-1) & MULT_11_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(0,0)<=signed(MULT_11_5(0,0)(MULT_SIZE-1) & MULT_11_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(0,0)(MULT_SIZE-1) & MULT_11_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(0,0)<=signed(MULT_12_1(0,0)(MULT_SIZE-1) & MULT_12_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(0,0)(MULT_SIZE-1) & MULT_12_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(0,0)<=signed(MULT_12_3(0,0)(MULT_SIZE-1) & MULT_12_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(0,0)(MULT_SIZE-1) & MULT_12_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(0,0)<=signed(MULT_12_5(0,0)(MULT_SIZE-1) & MULT_12_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(0,0)(MULT_SIZE-1) & MULT_12_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(0,0)<=signed(MULT_13_1(0,0)(MULT_SIZE-1) & MULT_13_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(0,0)(MULT_SIZE-1) & MULT_13_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(0,0)<=signed(MULT_13_3(0,0)(MULT_SIZE-1) & MULT_13_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(0,0)(MULT_SIZE-1) & MULT_13_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(0,0)<=signed(MULT_13_5(0,0)(MULT_SIZE-1) & MULT_13_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(0,0)(MULT_SIZE-1) & MULT_13_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(0,0)<=signed(MULT_14_1(0,0)(MULT_SIZE-1) & MULT_14_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(0,0)(MULT_SIZE-1) & MULT_14_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(0,0)<=signed(MULT_14_3(0,0)(MULT_SIZE-1) & MULT_14_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(0,0)(MULT_SIZE-1) & MULT_14_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(0,0)<=signed(MULT_14_5(0,0)(MULT_SIZE-1) & MULT_14_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(0,0)(MULT_SIZE-1) & MULT_14_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(0,0)<=signed(MULT_15_1(0,0)(MULT_SIZE-1) & MULT_15_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(0,0)(MULT_SIZE-1) & MULT_15_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(0,0)<=signed(MULT_15_3(0,0)(MULT_SIZE-1) & MULT_15_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(0,0)(MULT_SIZE-1) & MULT_15_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(0,0)<=signed(MULT_15_5(0,0)(MULT_SIZE-1) & MULT_15_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(0,0)(MULT_SIZE-1) & MULT_15_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(0,0)<=signed(MULT_16_1(0,0)(MULT_SIZE-1) & MULT_16_1(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(0,0)(MULT_SIZE-1) & MULT_16_2(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(0,0)<=signed(MULT_16_3(0,0)(MULT_SIZE-1) & MULT_16_3(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(0,0)(MULT_SIZE-1) & MULT_16_4(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(0,0)<=signed(MULT_16_5(0,0)(MULT_SIZE-1) & MULT_16_5(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(0,0)(MULT_SIZE-1) & MULT_16_6(0,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(0,0) ------------------

			MULTS_1_1_1(0,1)<=signed(MULT_1_1(0,1)(MULT_SIZE-1) & MULT_1_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(0,1)(MULT_SIZE-1) & MULT_1_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(0,1)<=signed(MULT_1_3(0,1)(MULT_SIZE-1) & MULT_1_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(0,1)(MULT_SIZE-1) & MULT_1_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(0,1)<=signed(MULT_1_5(0,1)(MULT_SIZE-1) & MULT_1_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(0,1)(MULT_SIZE-1) & MULT_1_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(0,1)<=signed(MULT_2_1(0,1)(MULT_SIZE-1) & MULT_2_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(0,1)(MULT_SIZE-1) & MULT_2_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(0,1)<=signed(MULT_2_3(0,1)(MULT_SIZE-1) & MULT_2_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(0,1)(MULT_SIZE-1) & MULT_2_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(0,1)<=signed(MULT_2_5(0,1)(MULT_SIZE-1) & MULT_2_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(0,1)(MULT_SIZE-1) & MULT_2_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(0,1)<=signed(MULT_3_1(0,1)(MULT_SIZE-1) & MULT_3_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(0,1)(MULT_SIZE-1) & MULT_3_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(0,1)<=signed(MULT_3_3(0,1)(MULT_SIZE-1) & MULT_3_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(0,1)(MULT_SIZE-1) & MULT_3_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(0,1)<=signed(MULT_3_5(0,1)(MULT_SIZE-1) & MULT_3_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(0,1)(MULT_SIZE-1) & MULT_3_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(0,1)<=signed(MULT_4_1(0,1)(MULT_SIZE-1) & MULT_4_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(0,1)(MULT_SIZE-1) & MULT_4_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(0,1)<=signed(MULT_4_3(0,1)(MULT_SIZE-1) & MULT_4_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(0,1)(MULT_SIZE-1) & MULT_4_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(0,1)<=signed(MULT_4_5(0,1)(MULT_SIZE-1) & MULT_4_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(0,1)(MULT_SIZE-1) & MULT_4_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(0,1)<=signed(MULT_5_1(0,1)(MULT_SIZE-1) & MULT_5_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(0,1)(MULT_SIZE-1) & MULT_5_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(0,1)<=signed(MULT_5_3(0,1)(MULT_SIZE-1) & MULT_5_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(0,1)(MULT_SIZE-1) & MULT_5_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(0,1)<=signed(MULT_5_5(0,1)(MULT_SIZE-1) & MULT_5_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(0,1)(MULT_SIZE-1) & MULT_5_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(0,1)<=signed(MULT_6_1(0,1)(MULT_SIZE-1) & MULT_6_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(0,1)(MULT_SIZE-1) & MULT_6_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(0,1)<=signed(MULT_6_3(0,1)(MULT_SIZE-1) & MULT_6_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(0,1)(MULT_SIZE-1) & MULT_6_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(0,1)<=signed(MULT_6_5(0,1)(MULT_SIZE-1) & MULT_6_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(0,1)(MULT_SIZE-1) & MULT_6_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(0,1)<=signed(MULT_7_1(0,1)(MULT_SIZE-1) & MULT_7_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(0,1)(MULT_SIZE-1) & MULT_7_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(0,1)<=signed(MULT_7_3(0,1)(MULT_SIZE-1) & MULT_7_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(0,1)(MULT_SIZE-1) & MULT_7_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(0,1)<=signed(MULT_7_5(0,1)(MULT_SIZE-1) & MULT_7_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(0,1)(MULT_SIZE-1) & MULT_7_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(0,1)<=signed(MULT_8_1(0,1)(MULT_SIZE-1) & MULT_8_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(0,1)(MULT_SIZE-1) & MULT_8_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(0,1)<=signed(MULT_8_3(0,1)(MULT_SIZE-1) & MULT_8_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(0,1)(MULT_SIZE-1) & MULT_8_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(0,1)<=signed(MULT_8_5(0,1)(MULT_SIZE-1) & MULT_8_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(0,1)(MULT_SIZE-1) & MULT_8_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(0,1)<=signed(MULT_9_1(0,1)(MULT_SIZE-1) & MULT_9_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(0,1)(MULT_SIZE-1) & MULT_9_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(0,1)<=signed(MULT_9_3(0,1)(MULT_SIZE-1) & MULT_9_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(0,1)(MULT_SIZE-1) & MULT_9_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(0,1)<=signed(MULT_9_5(0,1)(MULT_SIZE-1) & MULT_9_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(0,1)(MULT_SIZE-1) & MULT_9_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(0,1)<=signed(MULT_10_1(0,1)(MULT_SIZE-1) & MULT_10_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(0,1)(MULT_SIZE-1) & MULT_10_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(0,1)<=signed(MULT_10_3(0,1)(MULT_SIZE-1) & MULT_10_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(0,1)(MULT_SIZE-1) & MULT_10_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(0,1)<=signed(MULT_10_5(0,1)(MULT_SIZE-1) & MULT_10_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(0,1)(MULT_SIZE-1) & MULT_10_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(0,1)<=signed(MULT_11_1(0,1)(MULT_SIZE-1) & MULT_11_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(0,1)(MULT_SIZE-1) & MULT_11_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(0,1)<=signed(MULT_11_3(0,1)(MULT_SIZE-1) & MULT_11_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(0,1)(MULT_SIZE-1) & MULT_11_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(0,1)<=signed(MULT_11_5(0,1)(MULT_SIZE-1) & MULT_11_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(0,1)(MULT_SIZE-1) & MULT_11_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(0,1)<=signed(MULT_12_1(0,1)(MULT_SIZE-1) & MULT_12_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(0,1)(MULT_SIZE-1) & MULT_12_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(0,1)<=signed(MULT_12_3(0,1)(MULT_SIZE-1) & MULT_12_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(0,1)(MULT_SIZE-1) & MULT_12_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(0,1)<=signed(MULT_12_5(0,1)(MULT_SIZE-1) & MULT_12_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(0,1)(MULT_SIZE-1) & MULT_12_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(0,1)<=signed(MULT_13_1(0,1)(MULT_SIZE-1) & MULT_13_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(0,1)(MULT_SIZE-1) & MULT_13_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(0,1)<=signed(MULT_13_3(0,1)(MULT_SIZE-1) & MULT_13_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(0,1)(MULT_SIZE-1) & MULT_13_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(0,1)<=signed(MULT_13_5(0,1)(MULT_SIZE-1) & MULT_13_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(0,1)(MULT_SIZE-1) & MULT_13_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(0,1)<=signed(MULT_14_1(0,1)(MULT_SIZE-1) & MULT_14_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(0,1)(MULT_SIZE-1) & MULT_14_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(0,1)<=signed(MULT_14_3(0,1)(MULT_SIZE-1) & MULT_14_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(0,1)(MULT_SIZE-1) & MULT_14_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(0,1)<=signed(MULT_14_5(0,1)(MULT_SIZE-1) & MULT_14_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(0,1)(MULT_SIZE-1) & MULT_14_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(0,1)<=signed(MULT_15_1(0,1)(MULT_SIZE-1) & MULT_15_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(0,1)(MULT_SIZE-1) & MULT_15_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(0,1)<=signed(MULT_15_3(0,1)(MULT_SIZE-1) & MULT_15_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(0,1)(MULT_SIZE-1) & MULT_15_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(0,1)<=signed(MULT_15_5(0,1)(MULT_SIZE-1) & MULT_15_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(0,1)(MULT_SIZE-1) & MULT_15_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(0,1)<=signed(MULT_16_1(0,1)(MULT_SIZE-1) & MULT_16_1(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(0,1)(MULT_SIZE-1) & MULT_16_2(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(0,1)<=signed(MULT_16_3(0,1)(MULT_SIZE-1) & MULT_16_3(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(0,1)(MULT_SIZE-1) & MULT_16_4(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(0,1)<=signed(MULT_16_5(0,1)(MULT_SIZE-1) & MULT_16_5(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(0,1)(MULT_SIZE-1) & MULT_16_6(0,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(0,1) ------------------

			MULTS_1_1_1(0,2)<=signed(MULT_1_1(0,2)(MULT_SIZE-1) & MULT_1_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(0,2)(MULT_SIZE-1) & MULT_1_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(0,2)<=signed(MULT_1_3(0,2)(MULT_SIZE-1) & MULT_1_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(0,2)(MULT_SIZE-1) & MULT_1_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(0,2)<=signed(MULT_1_5(0,2)(MULT_SIZE-1) & MULT_1_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(0,2)(MULT_SIZE-1) & MULT_1_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(0,2)<=signed(MULT_2_1(0,2)(MULT_SIZE-1) & MULT_2_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(0,2)(MULT_SIZE-1) & MULT_2_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(0,2)<=signed(MULT_2_3(0,2)(MULT_SIZE-1) & MULT_2_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(0,2)(MULT_SIZE-1) & MULT_2_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(0,2)<=signed(MULT_2_5(0,2)(MULT_SIZE-1) & MULT_2_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(0,2)(MULT_SIZE-1) & MULT_2_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(0,2)<=signed(MULT_3_1(0,2)(MULT_SIZE-1) & MULT_3_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(0,2)(MULT_SIZE-1) & MULT_3_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(0,2)<=signed(MULT_3_3(0,2)(MULT_SIZE-1) & MULT_3_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(0,2)(MULT_SIZE-1) & MULT_3_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(0,2)<=signed(MULT_3_5(0,2)(MULT_SIZE-1) & MULT_3_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(0,2)(MULT_SIZE-1) & MULT_3_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(0,2)<=signed(MULT_4_1(0,2)(MULT_SIZE-1) & MULT_4_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(0,2)(MULT_SIZE-1) & MULT_4_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(0,2)<=signed(MULT_4_3(0,2)(MULT_SIZE-1) & MULT_4_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(0,2)(MULT_SIZE-1) & MULT_4_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(0,2)<=signed(MULT_4_5(0,2)(MULT_SIZE-1) & MULT_4_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(0,2)(MULT_SIZE-1) & MULT_4_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(0,2)<=signed(MULT_5_1(0,2)(MULT_SIZE-1) & MULT_5_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(0,2)(MULT_SIZE-1) & MULT_5_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(0,2)<=signed(MULT_5_3(0,2)(MULT_SIZE-1) & MULT_5_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(0,2)(MULT_SIZE-1) & MULT_5_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(0,2)<=signed(MULT_5_5(0,2)(MULT_SIZE-1) & MULT_5_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(0,2)(MULT_SIZE-1) & MULT_5_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(0,2)<=signed(MULT_6_1(0,2)(MULT_SIZE-1) & MULT_6_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(0,2)(MULT_SIZE-1) & MULT_6_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(0,2)<=signed(MULT_6_3(0,2)(MULT_SIZE-1) & MULT_6_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(0,2)(MULT_SIZE-1) & MULT_6_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(0,2)<=signed(MULT_6_5(0,2)(MULT_SIZE-1) & MULT_6_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(0,2)(MULT_SIZE-1) & MULT_6_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(0,2)<=signed(MULT_7_1(0,2)(MULT_SIZE-1) & MULT_7_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(0,2)(MULT_SIZE-1) & MULT_7_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(0,2)<=signed(MULT_7_3(0,2)(MULT_SIZE-1) & MULT_7_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(0,2)(MULT_SIZE-1) & MULT_7_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(0,2)<=signed(MULT_7_5(0,2)(MULT_SIZE-1) & MULT_7_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(0,2)(MULT_SIZE-1) & MULT_7_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(0,2)<=signed(MULT_8_1(0,2)(MULT_SIZE-1) & MULT_8_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(0,2)(MULT_SIZE-1) & MULT_8_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(0,2)<=signed(MULT_8_3(0,2)(MULT_SIZE-1) & MULT_8_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(0,2)(MULT_SIZE-1) & MULT_8_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(0,2)<=signed(MULT_8_5(0,2)(MULT_SIZE-1) & MULT_8_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(0,2)(MULT_SIZE-1) & MULT_8_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(0,2)<=signed(MULT_9_1(0,2)(MULT_SIZE-1) & MULT_9_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(0,2)(MULT_SIZE-1) & MULT_9_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(0,2)<=signed(MULT_9_3(0,2)(MULT_SIZE-1) & MULT_9_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(0,2)(MULT_SIZE-1) & MULT_9_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(0,2)<=signed(MULT_9_5(0,2)(MULT_SIZE-1) & MULT_9_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(0,2)(MULT_SIZE-1) & MULT_9_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(0,2)<=signed(MULT_10_1(0,2)(MULT_SIZE-1) & MULT_10_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(0,2)(MULT_SIZE-1) & MULT_10_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(0,2)<=signed(MULT_10_3(0,2)(MULT_SIZE-1) & MULT_10_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(0,2)(MULT_SIZE-1) & MULT_10_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(0,2)<=signed(MULT_10_5(0,2)(MULT_SIZE-1) & MULT_10_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(0,2)(MULT_SIZE-1) & MULT_10_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(0,2)<=signed(MULT_11_1(0,2)(MULT_SIZE-1) & MULT_11_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(0,2)(MULT_SIZE-1) & MULT_11_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(0,2)<=signed(MULT_11_3(0,2)(MULT_SIZE-1) & MULT_11_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(0,2)(MULT_SIZE-1) & MULT_11_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(0,2)<=signed(MULT_11_5(0,2)(MULT_SIZE-1) & MULT_11_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(0,2)(MULT_SIZE-1) & MULT_11_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(0,2)<=signed(MULT_12_1(0,2)(MULT_SIZE-1) & MULT_12_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(0,2)(MULT_SIZE-1) & MULT_12_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(0,2)<=signed(MULT_12_3(0,2)(MULT_SIZE-1) & MULT_12_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(0,2)(MULT_SIZE-1) & MULT_12_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(0,2)<=signed(MULT_12_5(0,2)(MULT_SIZE-1) & MULT_12_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(0,2)(MULT_SIZE-1) & MULT_12_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(0,2)<=signed(MULT_13_1(0,2)(MULT_SIZE-1) & MULT_13_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(0,2)(MULT_SIZE-1) & MULT_13_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(0,2)<=signed(MULT_13_3(0,2)(MULT_SIZE-1) & MULT_13_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(0,2)(MULT_SIZE-1) & MULT_13_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(0,2)<=signed(MULT_13_5(0,2)(MULT_SIZE-1) & MULT_13_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(0,2)(MULT_SIZE-1) & MULT_13_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(0,2)<=signed(MULT_14_1(0,2)(MULT_SIZE-1) & MULT_14_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(0,2)(MULT_SIZE-1) & MULT_14_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(0,2)<=signed(MULT_14_3(0,2)(MULT_SIZE-1) & MULT_14_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(0,2)(MULT_SIZE-1) & MULT_14_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(0,2)<=signed(MULT_14_5(0,2)(MULT_SIZE-1) & MULT_14_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(0,2)(MULT_SIZE-1) & MULT_14_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(0,2)<=signed(MULT_15_1(0,2)(MULT_SIZE-1) & MULT_15_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(0,2)(MULT_SIZE-1) & MULT_15_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(0,2)<=signed(MULT_15_3(0,2)(MULT_SIZE-1) & MULT_15_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(0,2)(MULT_SIZE-1) & MULT_15_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(0,2)<=signed(MULT_15_5(0,2)(MULT_SIZE-1) & MULT_15_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(0,2)(MULT_SIZE-1) & MULT_15_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(0,2)<=signed(MULT_16_1(0,2)(MULT_SIZE-1) & MULT_16_1(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(0,2)(MULT_SIZE-1) & MULT_16_2(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(0,2)<=signed(MULT_16_3(0,2)(MULT_SIZE-1) & MULT_16_3(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(0,2)(MULT_SIZE-1) & MULT_16_4(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(0,2)<=signed(MULT_16_5(0,2)(MULT_SIZE-1) & MULT_16_5(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(0,2)(MULT_SIZE-1) & MULT_16_6(0,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(0,2) ------------------

			MULTS_1_1_1(0,3)<=signed(MULT_1_1(0,3)(MULT_SIZE-1) & MULT_1_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(0,3)(MULT_SIZE-1) & MULT_1_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(0,3)<=signed(MULT_1_3(0,3)(MULT_SIZE-1) & MULT_1_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(0,3)(MULT_SIZE-1) & MULT_1_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(0,3)<=signed(MULT_1_5(0,3)(MULT_SIZE-1) & MULT_1_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(0,3)(MULT_SIZE-1) & MULT_1_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(0,3)<=signed(MULT_2_1(0,3)(MULT_SIZE-1) & MULT_2_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(0,3)(MULT_SIZE-1) & MULT_2_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(0,3)<=signed(MULT_2_3(0,3)(MULT_SIZE-1) & MULT_2_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(0,3)(MULT_SIZE-1) & MULT_2_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(0,3)<=signed(MULT_2_5(0,3)(MULT_SIZE-1) & MULT_2_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(0,3)(MULT_SIZE-1) & MULT_2_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(0,3)<=signed(MULT_3_1(0,3)(MULT_SIZE-1) & MULT_3_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(0,3)(MULT_SIZE-1) & MULT_3_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(0,3)<=signed(MULT_3_3(0,3)(MULT_SIZE-1) & MULT_3_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(0,3)(MULT_SIZE-1) & MULT_3_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(0,3)<=signed(MULT_3_5(0,3)(MULT_SIZE-1) & MULT_3_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(0,3)(MULT_SIZE-1) & MULT_3_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(0,3)<=signed(MULT_4_1(0,3)(MULT_SIZE-1) & MULT_4_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(0,3)(MULT_SIZE-1) & MULT_4_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(0,3)<=signed(MULT_4_3(0,3)(MULT_SIZE-1) & MULT_4_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(0,3)(MULT_SIZE-1) & MULT_4_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(0,3)<=signed(MULT_4_5(0,3)(MULT_SIZE-1) & MULT_4_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(0,3)(MULT_SIZE-1) & MULT_4_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(0,3)<=signed(MULT_5_1(0,3)(MULT_SIZE-1) & MULT_5_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(0,3)(MULT_SIZE-1) & MULT_5_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(0,3)<=signed(MULT_5_3(0,3)(MULT_SIZE-1) & MULT_5_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(0,3)(MULT_SIZE-1) & MULT_5_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(0,3)<=signed(MULT_5_5(0,3)(MULT_SIZE-1) & MULT_5_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(0,3)(MULT_SIZE-1) & MULT_5_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(0,3)<=signed(MULT_6_1(0,3)(MULT_SIZE-1) & MULT_6_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(0,3)(MULT_SIZE-1) & MULT_6_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(0,3)<=signed(MULT_6_3(0,3)(MULT_SIZE-1) & MULT_6_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(0,3)(MULT_SIZE-1) & MULT_6_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(0,3)<=signed(MULT_6_5(0,3)(MULT_SIZE-1) & MULT_6_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(0,3)(MULT_SIZE-1) & MULT_6_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(0,3)<=signed(MULT_7_1(0,3)(MULT_SIZE-1) & MULT_7_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(0,3)(MULT_SIZE-1) & MULT_7_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(0,3)<=signed(MULT_7_3(0,3)(MULT_SIZE-1) & MULT_7_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(0,3)(MULT_SIZE-1) & MULT_7_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(0,3)<=signed(MULT_7_5(0,3)(MULT_SIZE-1) & MULT_7_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(0,3)(MULT_SIZE-1) & MULT_7_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(0,3)<=signed(MULT_8_1(0,3)(MULT_SIZE-1) & MULT_8_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(0,3)(MULT_SIZE-1) & MULT_8_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(0,3)<=signed(MULT_8_3(0,3)(MULT_SIZE-1) & MULT_8_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(0,3)(MULT_SIZE-1) & MULT_8_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(0,3)<=signed(MULT_8_5(0,3)(MULT_SIZE-1) & MULT_8_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(0,3)(MULT_SIZE-1) & MULT_8_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(0,3)<=signed(MULT_9_1(0,3)(MULT_SIZE-1) & MULT_9_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(0,3)(MULT_SIZE-1) & MULT_9_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(0,3)<=signed(MULT_9_3(0,3)(MULT_SIZE-1) & MULT_9_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(0,3)(MULT_SIZE-1) & MULT_9_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(0,3)<=signed(MULT_9_5(0,3)(MULT_SIZE-1) & MULT_9_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(0,3)(MULT_SIZE-1) & MULT_9_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(0,3)<=signed(MULT_10_1(0,3)(MULT_SIZE-1) & MULT_10_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(0,3)(MULT_SIZE-1) & MULT_10_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(0,3)<=signed(MULT_10_3(0,3)(MULT_SIZE-1) & MULT_10_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(0,3)(MULT_SIZE-1) & MULT_10_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(0,3)<=signed(MULT_10_5(0,3)(MULT_SIZE-1) & MULT_10_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(0,3)(MULT_SIZE-1) & MULT_10_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(0,3)<=signed(MULT_11_1(0,3)(MULT_SIZE-1) & MULT_11_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(0,3)(MULT_SIZE-1) & MULT_11_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(0,3)<=signed(MULT_11_3(0,3)(MULT_SIZE-1) & MULT_11_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(0,3)(MULT_SIZE-1) & MULT_11_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(0,3)<=signed(MULT_11_5(0,3)(MULT_SIZE-1) & MULT_11_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(0,3)(MULT_SIZE-1) & MULT_11_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(0,3)<=signed(MULT_12_1(0,3)(MULT_SIZE-1) & MULT_12_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(0,3)(MULT_SIZE-1) & MULT_12_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(0,3)<=signed(MULT_12_3(0,3)(MULT_SIZE-1) & MULT_12_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(0,3)(MULT_SIZE-1) & MULT_12_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(0,3)<=signed(MULT_12_5(0,3)(MULT_SIZE-1) & MULT_12_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(0,3)(MULT_SIZE-1) & MULT_12_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(0,3)<=signed(MULT_13_1(0,3)(MULT_SIZE-1) & MULT_13_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(0,3)(MULT_SIZE-1) & MULT_13_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(0,3)<=signed(MULT_13_3(0,3)(MULT_SIZE-1) & MULT_13_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(0,3)(MULT_SIZE-1) & MULT_13_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(0,3)<=signed(MULT_13_5(0,3)(MULT_SIZE-1) & MULT_13_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(0,3)(MULT_SIZE-1) & MULT_13_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(0,3)<=signed(MULT_14_1(0,3)(MULT_SIZE-1) & MULT_14_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(0,3)(MULT_SIZE-1) & MULT_14_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(0,3)<=signed(MULT_14_3(0,3)(MULT_SIZE-1) & MULT_14_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(0,3)(MULT_SIZE-1) & MULT_14_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(0,3)<=signed(MULT_14_5(0,3)(MULT_SIZE-1) & MULT_14_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(0,3)(MULT_SIZE-1) & MULT_14_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(0,3)<=signed(MULT_15_1(0,3)(MULT_SIZE-1) & MULT_15_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(0,3)(MULT_SIZE-1) & MULT_15_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(0,3)<=signed(MULT_15_3(0,3)(MULT_SIZE-1) & MULT_15_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(0,3)(MULT_SIZE-1) & MULT_15_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(0,3)<=signed(MULT_15_5(0,3)(MULT_SIZE-1) & MULT_15_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(0,3)(MULT_SIZE-1) & MULT_15_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(0,3)<=signed(MULT_16_1(0,3)(MULT_SIZE-1) & MULT_16_1(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(0,3)(MULT_SIZE-1) & MULT_16_2(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(0,3)<=signed(MULT_16_3(0,3)(MULT_SIZE-1) & MULT_16_3(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(0,3)(MULT_SIZE-1) & MULT_16_4(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(0,3)<=signed(MULT_16_5(0,3)(MULT_SIZE-1) & MULT_16_5(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(0,3)(MULT_SIZE-1) & MULT_16_6(0,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(0,3) ------------------

			MULTS_1_1_1(0,4)<=signed(MULT_1_1(0,4)(MULT_SIZE-1) & MULT_1_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(0,4)(MULT_SIZE-1) & MULT_1_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(0,4)<=signed(MULT_1_3(0,4)(MULT_SIZE-1) & MULT_1_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(0,4)(MULT_SIZE-1) & MULT_1_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(0,4)<=signed(MULT_1_5(0,4)(MULT_SIZE-1) & MULT_1_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(0,4)(MULT_SIZE-1) & MULT_1_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(0,4)<=signed(MULT_2_1(0,4)(MULT_SIZE-1) & MULT_2_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(0,4)(MULT_SIZE-1) & MULT_2_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(0,4)<=signed(MULT_2_3(0,4)(MULT_SIZE-1) & MULT_2_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(0,4)(MULT_SIZE-1) & MULT_2_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(0,4)<=signed(MULT_2_5(0,4)(MULT_SIZE-1) & MULT_2_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(0,4)(MULT_SIZE-1) & MULT_2_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(0,4)<=signed(MULT_3_1(0,4)(MULT_SIZE-1) & MULT_3_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(0,4)(MULT_SIZE-1) & MULT_3_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(0,4)<=signed(MULT_3_3(0,4)(MULT_SIZE-1) & MULT_3_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(0,4)(MULT_SIZE-1) & MULT_3_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(0,4)<=signed(MULT_3_5(0,4)(MULT_SIZE-1) & MULT_3_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(0,4)(MULT_SIZE-1) & MULT_3_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(0,4)<=signed(MULT_4_1(0,4)(MULT_SIZE-1) & MULT_4_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(0,4)(MULT_SIZE-1) & MULT_4_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(0,4)<=signed(MULT_4_3(0,4)(MULT_SIZE-1) & MULT_4_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(0,4)(MULT_SIZE-1) & MULT_4_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(0,4)<=signed(MULT_4_5(0,4)(MULT_SIZE-1) & MULT_4_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(0,4)(MULT_SIZE-1) & MULT_4_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(0,4)<=signed(MULT_5_1(0,4)(MULT_SIZE-1) & MULT_5_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(0,4)(MULT_SIZE-1) & MULT_5_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(0,4)<=signed(MULT_5_3(0,4)(MULT_SIZE-1) & MULT_5_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(0,4)(MULT_SIZE-1) & MULT_5_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(0,4)<=signed(MULT_5_5(0,4)(MULT_SIZE-1) & MULT_5_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(0,4)(MULT_SIZE-1) & MULT_5_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(0,4)<=signed(MULT_6_1(0,4)(MULT_SIZE-1) & MULT_6_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(0,4)(MULT_SIZE-1) & MULT_6_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(0,4)<=signed(MULT_6_3(0,4)(MULT_SIZE-1) & MULT_6_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(0,4)(MULT_SIZE-1) & MULT_6_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(0,4)<=signed(MULT_6_5(0,4)(MULT_SIZE-1) & MULT_6_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(0,4)(MULT_SIZE-1) & MULT_6_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(0,4)<=signed(MULT_7_1(0,4)(MULT_SIZE-1) & MULT_7_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(0,4)(MULT_SIZE-1) & MULT_7_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(0,4)<=signed(MULT_7_3(0,4)(MULT_SIZE-1) & MULT_7_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(0,4)(MULT_SIZE-1) & MULT_7_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(0,4)<=signed(MULT_7_5(0,4)(MULT_SIZE-1) & MULT_7_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(0,4)(MULT_SIZE-1) & MULT_7_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(0,4)<=signed(MULT_8_1(0,4)(MULT_SIZE-1) & MULT_8_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(0,4)(MULT_SIZE-1) & MULT_8_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(0,4)<=signed(MULT_8_3(0,4)(MULT_SIZE-1) & MULT_8_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(0,4)(MULT_SIZE-1) & MULT_8_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(0,4)<=signed(MULT_8_5(0,4)(MULT_SIZE-1) & MULT_8_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(0,4)(MULT_SIZE-1) & MULT_8_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(0,4)<=signed(MULT_9_1(0,4)(MULT_SIZE-1) & MULT_9_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(0,4)(MULT_SIZE-1) & MULT_9_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(0,4)<=signed(MULT_9_3(0,4)(MULT_SIZE-1) & MULT_9_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(0,4)(MULT_SIZE-1) & MULT_9_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(0,4)<=signed(MULT_9_5(0,4)(MULT_SIZE-1) & MULT_9_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(0,4)(MULT_SIZE-1) & MULT_9_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(0,4)<=signed(MULT_10_1(0,4)(MULT_SIZE-1) & MULT_10_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(0,4)(MULT_SIZE-1) & MULT_10_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(0,4)<=signed(MULT_10_3(0,4)(MULT_SIZE-1) & MULT_10_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(0,4)(MULT_SIZE-1) & MULT_10_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(0,4)<=signed(MULT_10_5(0,4)(MULT_SIZE-1) & MULT_10_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(0,4)(MULT_SIZE-1) & MULT_10_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(0,4)<=signed(MULT_11_1(0,4)(MULT_SIZE-1) & MULT_11_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(0,4)(MULT_SIZE-1) & MULT_11_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(0,4)<=signed(MULT_11_3(0,4)(MULT_SIZE-1) & MULT_11_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(0,4)(MULT_SIZE-1) & MULT_11_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(0,4)<=signed(MULT_11_5(0,4)(MULT_SIZE-1) & MULT_11_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(0,4)(MULT_SIZE-1) & MULT_11_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(0,4)<=signed(MULT_12_1(0,4)(MULT_SIZE-1) & MULT_12_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(0,4)(MULT_SIZE-1) & MULT_12_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(0,4)<=signed(MULT_12_3(0,4)(MULT_SIZE-1) & MULT_12_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(0,4)(MULT_SIZE-1) & MULT_12_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(0,4)<=signed(MULT_12_5(0,4)(MULT_SIZE-1) & MULT_12_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(0,4)(MULT_SIZE-1) & MULT_12_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(0,4)<=signed(MULT_13_1(0,4)(MULT_SIZE-1) & MULT_13_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(0,4)(MULT_SIZE-1) & MULT_13_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(0,4)<=signed(MULT_13_3(0,4)(MULT_SIZE-1) & MULT_13_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(0,4)(MULT_SIZE-1) & MULT_13_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(0,4)<=signed(MULT_13_5(0,4)(MULT_SIZE-1) & MULT_13_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(0,4)(MULT_SIZE-1) & MULT_13_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(0,4)<=signed(MULT_14_1(0,4)(MULT_SIZE-1) & MULT_14_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(0,4)(MULT_SIZE-1) & MULT_14_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(0,4)<=signed(MULT_14_3(0,4)(MULT_SIZE-1) & MULT_14_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(0,4)(MULT_SIZE-1) & MULT_14_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(0,4)<=signed(MULT_14_5(0,4)(MULT_SIZE-1) & MULT_14_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(0,4)(MULT_SIZE-1) & MULT_14_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(0,4)<=signed(MULT_15_1(0,4)(MULT_SIZE-1) & MULT_15_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(0,4)(MULT_SIZE-1) & MULT_15_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(0,4)<=signed(MULT_15_3(0,4)(MULT_SIZE-1) & MULT_15_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(0,4)(MULT_SIZE-1) & MULT_15_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(0,4)<=signed(MULT_15_5(0,4)(MULT_SIZE-1) & MULT_15_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(0,4)(MULT_SIZE-1) & MULT_15_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(0,4)<=signed(MULT_16_1(0,4)(MULT_SIZE-1) & MULT_16_1(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(0,4)(MULT_SIZE-1) & MULT_16_2(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(0,4)<=signed(MULT_16_3(0,4)(MULT_SIZE-1) & MULT_16_3(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(0,4)(MULT_SIZE-1) & MULT_16_4(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(0,4)<=signed(MULT_16_5(0,4)(MULT_SIZE-1) & MULT_16_5(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(0,4)(MULT_SIZE-1) & MULT_16_6(0,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(0,4) ------------------

			MULTS_1_1_1(1,0)<=signed(MULT_1_1(1,0)(MULT_SIZE-1) & MULT_1_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(1,0)(MULT_SIZE-1) & MULT_1_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(1,0)<=signed(MULT_1_3(1,0)(MULT_SIZE-1) & MULT_1_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(1,0)(MULT_SIZE-1) & MULT_1_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(1,0)<=signed(MULT_1_5(1,0)(MULT_SIZE-1) & MULT_1_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(1,0)(MULT_SIZE-1) & MULT_1_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(1,0)<=signed(MULT_2_1(1,0)(MULT_SIZE-1) & MULT_2_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(1,0)(MULT_SIZE-1) & MULT_2_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(1,0)<=signed(MULT_2_3(1,0)(MULT_SIZE-1) & MULT_2_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(1,0)(MULT_SIZE-1) & MULT_2_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(1,0)<=signed(MULT_2_5(1,0)(MULT_SIZE-1) & MULT_2_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(1,0)(MULT_SIZE-1) & MULT_2_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(1,0)<=signed(MULT_3_1(1,0)(MULT_SIZE-1) & MULT_3_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(1,0)(MULT_SIZE-1) & MULT_3_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(1,0)<=signed(MULT_3_3(1,0)(MULT_SIZE-1) & MULT_3_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(1,0)(MULT_SIZE-1) & MULT_3_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(1,0)<=signed(MULT_3_5(1,0)(MULT_SIZE-1) & MULT_3_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(1,0)(MULT_SIZE-1) & MULT_3_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(1,0)<=signed(MULT_4_1(1,0)(MULT_SIZE-1) & MULT_4_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(1,0)(MULT_SIZE-1) & MULT_4_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(1,0)<=signed(MULT_4_3(1,0)(MULT_SIZE-1) & MULT_4_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(1,0)(MULT_SIZE-1) & MULT_4_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(1,0)<=signed(MULT_4_5(1,0)(MULT_SIZE-1) & MULT_4_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(1,0)(MULT_SIZE-1) & MULT_4_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(1,0)<=signed(MULT_5_1(1,0)(MULT_SIZE-1) & MULT_5_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(1,0)(MULT_SIZE-1) & MULT_5_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(1,0)<=signed(MULT_5_3(1,0)(MULT_SIZE-1) & MULT_5_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(1,0)(MULT_SIZE-1) & MULT_5_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(1,0)<=signed(MULT_5_5(1,0)(MULT_SIZE-1) & MULT_5_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(1,0)(MULT_SIZE-1) & MULT_5_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(1,0)<=signed(MULT_6_1(1,0)(MULT_SIZE-1) & MULT_6_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(1,0)(MULT_SIZE-1) & MULT_6_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(1,0)<=signed(MULT_6_3(1,0)(MULT_SIZE-1) & MULT_6_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(1,0)(MULT_SIZE-1) & MULT_6_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(1,0)<=signed(MULT_6_5(1,0)(MULT_SIZE-1) & MULT_6_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(1,0)(MULT_SIZE-1) & MULT_6_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(1,0)<=signed(MULT_7_1(1,0)(MULT_SIZE-1) & MULT_7_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(1,0)(MULT_SIZE-1) & MULT_7_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(1,0)<=signed(MULT_7_3(1,0)(MULT_SIZE-1) & MULT_7_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(1,0)(MULT_SIZE-1) & MULT_7_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(1,0)<=signed(MULT_7_5(1,0)(MULT_SIZE-1) & MULT_7_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(1,0)(MULT_SIZE-1) & MULT_7_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(1,0)<=signed(MULT_8_1(1,0)(MULT_SIZE-1) & MULT_8_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(1,0)(MULT_SIZE-1) & MULT_8_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(1,0)<=signed(MULT_8_3(1,0)(MULT_SIZE-1) & MULT_8_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(1,0)(MULT_SIZE-1) & MULT_8_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(1,0)<=signed(MULT_8_5(1,0)(MULT_SIZE-1) & MULT_8_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(1,0)(MULT_SIZE-1) & MULT_8_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(1,0)<=signed(MULT_9_1(1,0)(MULT_SIZE-1) & MULT_9_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(1,0)(MULT_SIZE-1) & MULT_9_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(1,0)<=signed(MULT_9_3(1,0)(MULT_SIZE-1) & MULT_9_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(1,0)(MULT_SIZE-1) & MULT_9_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(1,0)<=signed(MULT_9_5(1,0)(MULT_SIZE-1) & MULT_9_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(1,0)(MULT_SIZE-1) & MULT_9_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(1,0)<=signed(MULT_10_1(1,0)(MULT_SIZE-1) & MULT_10_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(1,0)(MULT_SIZE-1) & MULT_10_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(1,0)<=signed(MULT_10_3(1,0)(MULT_SIZE-1) & MULT_10_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(1,0)(MULT_SIZE-1) & MULT_10_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(1,0)<=signed(MULT_10_5(1,0)(MULT_SIZE-1) & MULT_10_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(1,0)(MULT_SIZE-1) & MULT_10_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(1,0)<=signed(MULT_11_1(1,0)(MULT_SIZE-1) & MULT_11_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(1,0)(MULT_SIZE-1) & MULT_11_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(1,0)<=signed(MULT_11_3(1,0)(MULT_SIZE-1) & MULT_11_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(1,0)(MULT_SIZE-1) & MULT_11_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(1,0)<=signed(MULT_11_5(1,0)(MULT_SIZE-1) & MULT_11_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(1,0)(MULT_SIZE-1) & MULT_11_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(1,0)<=signed(MULT_12_1(1,0)(MULT_SIZE-1) & MULT_12_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(1,0)(MULT_SIZE-1) & MULT_12_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(1,0)<=signed(MULT_12_3(1,0)(MULT_SIZE-1) & MULT_12_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(1,0)(MULT_SIZE-1) & MULT_12_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(1,0)<=signed(MULT_12_5(1,0)(MULT_SIZE-1) & MULT_12_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(1,0)(MULT_SIZE-1) & MULT_12_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(1,0)<=signed(MULT_13_1(1,0)(MULT_SIZE-1) & MULT_13_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(1,0)(MULT_SIZE-1) & MULT_13_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(1,0)<=signed(MULT_13_3(1,0)(MULT_SIZE-1) & MULT_13_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(1,0)(MULT_SIZE-1) & MULT_13_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(1,0)<=signed(MULT_13_5(1,0)(MULT_SIZE-1) & MULT_13_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(1,0)(MULT_SIZE-1) & MULT_13_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(1,0)<=signed(MULT_14_1(1,0)(MULT_SIZE-1) & MULT_14_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(1,0)(MULT_SIZE-1) & MULT_14_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(1,0)<=signed(MULT_14_3(1,0)(MULT_SIZE-1) & MULT_14_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(1,0)(MULT_SIZE-1) & MULT_14_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(1,0)<=signed(MULT_14_5(1,0)(MULT_SIZE-1) & MULT_14_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(1,0)(MULT_SIZE-1) & MULT_14_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(1,0)<=signed(MULT_15_1(1,0)(MULT_SIZE-1) & MULT_15_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(1,0)(MULT_SIZE-1) & MULT_15_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(1,0)<=signed(MULT_15_3(1,0)(MULT_SIZE-1) & MULT_15_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(1,0)(MULT_SIZE-1) & MULT_15_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(1,0)<=signed(MULT_15_5(1,0)(MULT_SIZE-1) & MULT_15_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(1,0)(MULT_SIZE-1) & MULT_15_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(1,0)<=signed(MULT_16_1(1,0)(MULT_SIZE-1) & MULT_16_1(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(1,0)(MULT_SIZE-1) & MULT_16_2(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(1,0)<=signed(MULT_16_3(1,0)(MULT_SIZE-1) & MULT_16_3(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(1,0)(MULT_SIZE-1) & MULT_16_4(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(1,0)<=signed(MULT_16_5(1,0)(MULT_SIZE-1) & MULT_16_5(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(1,0)(MULT_SIZE-1) & MULT_16_6(1,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(1,0) ------------------

			MULTS_1_1_1(1,1)<=signed(MULT_1_1(1,1)(MULT_SIZE-1) & MULT_1_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(1,1)(MULT_SIZE-1) & MULT_1_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(1,1)<=signed(MULT_1_3(1,1)(MULT_SIZE-1) & MULT_1_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(1,1)(MULT_SIZE-1) & MULT_1_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(1,1)<=signed(MULT_1_5(1,1)(MULT_SIZE-1) & MULT_1_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(1,1)(MULT_SIZE-1) & MULT_1_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(1,1)<=signed(MULT_2_1(1,1)(MULT_SIZE-1) & MULT_2_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(1,1)(MULT_SIZE-1) & MULT_2_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(1,1)<=signed(MULT_2_3(1,1)(MULT_SIZE-1) & MULT_2_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(1,1)(MULT_SIZE-1) & MULT_2_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(1,1)<=signed(MULT_2_5(1,1)(MULT_SIZE-1) & MULT_2_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(1,1)(MULT_SIZE-1) & MULT_2_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(1,1)<=signed(MULT_3_1(1,1)(MULT_SIZE-1) & MULT_3_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(1,1)(MULT_SIZE-1) & MULT_3_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(1,1)<=signed(MULT_3_3(1,1)(MULT_SIZE-1) & MULT_3_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(1,1)(MULT_SIZE-1) & MULT_3_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(1,1)<=signed(MULT_3_5(1,1)(MULT_SIZE-1) & MULT_3_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(1,1)(MULT_SIZE-1) & MULT_3_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(1,1)<=signed(MULT_4_1(1,1)(MULT_SIZE-1) & MULT_4_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(1,1)(MULT_SIZE-1) & MULT_4_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(1,1)<=signed(MULT_4_3(1,1)(MULT_SIZE-1) & MULT_4_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(1,1)(MULT_SIZE-1) & MULT_4_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(1,1)<=signed(MULT_4_5(1,1)(MULT_SIZE-1) & MULT_4_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(1,1)(MULT_SIZE-1) & MULT_4_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(1,1)<=signed(MULT_5_1(1,1)(MULT_SIZE-1) & MULT_5_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(1,1)(MULT_SIZE-1) & MULT_5_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(1,1)<=signed(MULT_5_3(1,1)(MULT_SIZE-1) & MULT_5_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(1,1)(MULT_SIZE-1) & MULT_5_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(1,1)<=signed(MULT_5_5(1,1)(MULT_SIZE-1) & MULT_5_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(1,1)(MULT_SIZE-1) & MULT_5_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(1,1)<=signed(MULT_6_1(1,1)(MULT_SIZE-1) & MULT_6_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(1,1)(MULT_SIZE-1) & MULT_6_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(1,1)<=signed(MULT_6_3(1,1)(MULT_SIZE-1) & MULT_6_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(1,1)(MULT_SIZE-1) & MULT_6_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(1,1)<=signed(MULT_6_5(1,1)(MULT_SIZE-1) & MULT_6_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(1,1)(MULT_SIZE-1) & MULT_6_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(1,1)<=signed(MULT_7_1(1,1)(MULT_SIZE-1) & MULT_7_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(1,1)(MULT_SIZE-1) & MULT_7_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(1,1)<=signed(MULT_7_3(1,1)(MULT_SIZE-1) & MULT_7_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(1,1)(MULT_SIZE-1) & MULT_7_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(1,1)<=signed(MULT_7_5(1,1)(MULT_SIZE-1) & MULT_7_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(1,1)(MULT_SIZE-1) & MULT_7_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(1,1)<=signed(MULT_8_1(1,1)(MULT_SIZE-1) & MULT_8_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(1,1)(MULT_SIZE-1) & MULT_8_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(1,1)<=signed(MULT_8_3(1,1)(MULT_SIZE-1) & MULT_8_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(1,1)(MULT_SIZE-1) & MULT_8_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(1,1)<=signed(MULT_8_5(1,1)(MULT_SIZE-1) & MULT_8_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(1,1)(MULT_SIZE-1) & MULT_8_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(1,1)<=signed(MULT_9_1(1,1)(MULT_SIZE-1) & MULT_9_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(1,1)(MULT_SIZE-1) & MULT_9_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(1,1)<=signed(MULT_9_3(1,1)(MULT_SIZE-1) & MULT_9_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(1,1)(MULT_SIZE-1) & MULT_9_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(1,1)<=signed(MULT_9_5(1,1)(MULT_SIZE-1) & MULT_9_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(1,1)(MULT_SIZE-1) & MULT_9_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(1,1)<=signed(MULT_10_1(1,1)(MULT_SIZE-1) & MULT_10_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(1,1)(MULT_SIZE-1) & MULT_10_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(1,1)<=signed(MULT_10_3(1,1)(MULT_SIZE-1) & MULT_10_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(1,1)(MULT_SIZE-1) & MULT_10_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(1,1)<=signed(MULT_10_5(1,1)(MULT_SIZE-1) & MULT_10_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(1,1)(MULT_SIZE-1) & MULT_10_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(1,1)<=signed(MULT_11_1(1,1)(MULT_SIZE-1) & MULT_11_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(1,1)(MULT_SIZE-1) & MULT_11_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(1,1)<=signed(MULT_11_3(1,1)(MULT_SIZE-1) & MULT_11_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(1,1)(MULT_SIZE-1) & MULT_11_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(1,1)<=signed(MULT_11_5(1,1)(MULT_SIZE-1) & MULT_11_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(1,1)(MULT_SIZE-1) & MULT_11_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(1,1)<=signed(MULT_12_1(1,1)(MULT_SIZE-1) & MULT_12_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(1,1)(MULT_SIZE-1) & MULT_12_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(1,1)<=signed(MULT_12_3(1,1)(MULT_SIZE-1) & MULT_12_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(1,1)(MULT_SIZE-1) & MULT_12_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(1,1)<=signed(MULT_12_5(1,1)(MULT_SIZE-1) & MULT_12_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(1,1)(MULT_SIZE-1) & MULT_12_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(1,1)<=signed(MULT_13_1(1,1)(MULT_SIZE-1) & MULT_13_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(1,1)(MULT_SIZE-1) & MULT_13_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(1,1)<=signed(MULT_13_3(1,1)(MULT_SIZE-1) & MULT_13_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(1,1)(MULT_SIZE-1) & MULT_13_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(1,1)<=signed(MULT_13_5(1,1)(MULT_SIZE-1) & MULT_13_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(1,1)(MULT_SIZE-1) & MULT_13_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(1,1)<=signed(MULT_14_1(1,1)(MULT_SIZE-1) & MULT_14_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(1,1)(MULT_SIZE-1) & MULT_14_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(1,1)<=signed(MULT_14_3(1,1)(MULT_SIZE-1) & MULT_14_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(1,1)(MULT_SIZE-1) & MULT_14_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(1,1)<=signed(MULT_14_5(1,1)(MULT_SIZE-1) & MULT_14_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(1,1)(MULT_SIZE-1) & MULT_14_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(1,1)<=signed(MULT_15_1(1,1)(MULT_SIZE-1) & MULT_15_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(1,1)(MULT_SIZE-1) & MULT_15_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(1,1)<=signed(MULT_15_3(1,1)(MULT_SIZE-1) & MULT_15_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(1,1)(MULT_SIZE-1) & MULT_15_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(1,1)<=signed(MULT_15_5(1,1)(MULT_SIZE-1) & MULT_15_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(1,1)(MULT_SIZE-1) & MULT_15_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(1,1)<=signed(MULT_16_1(1,1)(MULT_SIZE-1) & MULT_16_1(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(1,1)(MULT_SIZE-1) & MULT_16_2(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(1,1)<=signed(MULT_16_3(1,1)(MULT_SIZE-1) & MULT_16_3(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(1,1)(MULT_SIZE-1) & MULT_16_4(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(1,1)<=signed(MULT_16_5(1,1)(MULT_SIZE-1) & MULT_16_5(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(1,1)(MULT_SIZE-1) & MULT_16_6(1,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(1,1) ------------------

			MULTS_1_1_1(1,2)<=signed(MULT_1_1(1,2)(MULT_SIZE-1) & MULT_1_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(1,2)(MULT_SIZE-1) & MULT_1_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(1,2)<=signed(MULT_1_3(1,2)(MULT_SIZE-1) & MULT_1_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(1,2)(MULT_SIZE-1) & MULT_1_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(1,2)<=signed(MULT_1_5(1,2)(MULT_SIZE-1) & MULT_1_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(1,2)(MULT_SIZE-1) & MULT_1_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(1,2)<=signed(MULT_2_1(1,2)(MULT_SIZE-1) & MULT_2_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(1,2)(MULT_SIZE-1) & MULT_2_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(1,2)<=signed(MULT_2_3(1,2)(MULT_SIZE-1) & MULT_2_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(1,2)(MULT_SIZE-1) & MULT_2_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(1,2)<=signed(MULT_2_5(1,2)(MULT_SIZE-1) & MULT_2_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(1,2)(MULT_SIZE-1) & MULT_2_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(1,2)<=signed(MULT_3_1(1,2)(MULT_SIZE-1) & MULT_3_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(1,2)(MULT_SIZE-1) & MULT_3_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(1,2)<=signed(MULT_3_3(1,2)(MULT_SIZE-1) & MULT_3_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(1,2)(MULT_SIZE-1) & MULT_3_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(1,2)<=signed(MULT_3_5(1,2)(MULT_SIZE-1) & MULT_3_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(1,2)(MULT_SIZE-1) & MULT_3_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(1,2)<=signed(MULT_4_1(1,2)(MULT_SIZE-1) & MULT_4_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(1,2)(MULT_SIZE-1) & MULT_4_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(1,2)<=signed(MULT_4_3(1,2)(MULT_SIZE-1) & MULT_4_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(1,2)(MULT_SIZE-1) & MULT_4_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(1,2)<=signed(MULT_4_5(1,2)(MULT_SIZE-1) & MULT_4_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(1,2)(MULT_SIZE-1) & MULT_4_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(1,2)<=signed(MULT_5_1(1,2)(MULT_SIZE-1) & MULT_5_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(1,2)(MULT_SIZE-1) & MULT_5_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(1,2)<=signed(MULT_5_3(1,2)(MULT_SIZE-1) & MULT_5_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(1,2)(MULT_SIZE-1) & MULT_5_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(1,2)<=signed(MULT_5_5(1,2)(MULT_SIZE-1) & MULT_5_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(1,2)(MULT_SIZE-1) & MULT_5_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(1,2)<=signed(MULT_6_1(1,2)(MULT_SIZE-1) & MULT_6_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(1,2)(MULT_SIZE-1) & MULT_6_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(1,2)<=signed(MULT_6_3(1,2)(MULT_SIZE-1) & MULT_6_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(1,2)(MULT_SIZE-1) & MULT_6_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(1,2)<=signed(MULT_6_5(1,2)(MULT_SIZE-1) & MULT_6_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(1,2)(MULT_SIZE-1) & MULT_6_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(1,2)<=signed(MULT_7_1(1,2)(MULT_SIZE-1) & MULT_7_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(1,2)(MULT_SIZE-1) & MULT_7_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(1,2)<=signed(MULT_7_3(1,2)(MULT_SIZE-1) & MULT_7_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(1,2)(MULT_SIZE-1) & MULT_7_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(1,2)<=signed(MULT_7_5(1,2)(MULT_SIZE-1) & MULT_7_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(1,2)(MULT_SIZE-1) & MULT_7_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(1,2)<=signed(MULT_8_1(1,2)(MULT_SIZE-1) & MULT_8_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(1,2)(MULT_SIZE-1) & MULT_8_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(1,2)<=signed(MULT_8_3(1,2)(MULT_SIZE-1) & MULT_8_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(1,2)(MULT_SIZE-1) & MULT_8_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(1,2)<=signed(MULT_8_5(1,2)(MULT_SIZE-1) & MULT_8_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(1,2)(MULT_SIZE-1) & MULT_8_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(1,2)<=signed(MULT_9_1(1,2)(MULT_SIZE-1) & MULT_9_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(1,2)(MULT_SIZE-1) & MULT_9_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(1,2)<=signed(MULT_9_3(1,2)(MULT_SIZE-1) & MULT_9_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(1,2)(MULT_SIZE-1) & MULT_9_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(1,2)<=signed(MULT_9_5(1,2)(MULT_SIZE-1) & MULT_9_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(1,2)(MULT_SIZE-1) & MULT_9_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(1,2)<=signed(MULT_10_1(1,2)(MULT_SIZE-1) & MULT_10_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(1,2)(MULT_SIZE-1) & MULT_10_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(1,2)<=signed(MULT_10_3(1,2)(MULT_SIZE-1) & MULT_10_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(1,2)(MULT_SIZE-1) & MULT_10_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(1,2)<=signed(MULT_10_5(1,2)(MULT_SIZE-1) & MULT_10_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(1,2)(MULT_SIZE-1) & MULT_10_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(1,2)<=signed(MULT_11_1(1,2)(MULT_SIZE-1) & MULT_11_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(1,2)(MULT_SIZE-1) & MULT_11_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(1,2)<=signed(MULT_11_3(1,2)(MULT_SIZE-1) & MULT_11_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(1,2)(MULT_SIZE-1) & MULT_11_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(1,2)<=signed(MULT_11_5(1,2)(MULT_SIZE-1) & MULT_11_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(1,2)(MULT_SIZE-1) & MULT_11_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(1,2)<=signed(MULT_12_1(1,2)(MULT_SIZE-1) & MULT_12_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(1,2)(MULT_SIZE-1) & MULT_12_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(1,2)<=signed(MULT_12_3(1,2)(MULT_SIZE-1) & MULT_12_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(1,2)(MULT_SIZE-1) & MULT_12_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(1,2)<=signed(MULT_12_5(1,2)(MULT_SIZE-1) & MULT_12_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(1,2)(MULT_SIZE-1) & MULT_12_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(1,2)<=signed(MULT_13_1(1,2)(MULT_SIZE-1) & MULT_13_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(1,2)(MULT_SIZE-1) & MULT_13_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(1,2)<=signed(MULT_13_3(1,2)(MULT_SIZE-1) & MULT_13_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(1,2)(MULT_SIZE-1) & MULT_13_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(1,2)<=signed(MULT_13_5(1,2)(MULT_SIZE-1) & MULT_13_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(1,2)(MULT_SIZE-1) & MULT_13_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(1,2)<=signed(MULT_14_1(1,2)(MULT_SIZE-1) & MULT_14_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(1,2)(MULT_SIZE-1) & MULT_14_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(1,2)<=signed(MULT_14_3(1,2)(MULT_SIZE-1) & MULT_14_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(1,2)(MULT_SIZE-1) & MULT_14_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(1,2)<=signed(MULT_14_5(1,2)(MULT_SIZE-1) & MULT_14_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(1,2)(MULT_SIZE-1) & MULT_14_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(1,2)<=signed(MULT_15_1(1,2)(MULT_SIZE-1) & MULT_15_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(1,2)(MULT_SIZE-1) & MULT_15_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(1,2)<=signed(MULT_15_3(1,2)(MULT_SIZE-1) & MULT_15_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(1,2)(MULT_SIZE-1) & MULT_15_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(1,2)<=signed(MULT_15_5(1,2)(MULT_SIZE-1) & MULT_15_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(1,2)(MULT_SIZE-1) & MULT_15_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(1,2)<=signed(MULT_16_1(1,2)(MULT_SIZE-1) & MULT_16_1(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(1,2)(MULT_SIZE-1) & MULT_16_2(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(1,2)<=signed(MULT_16_3(1,2)(MULT_SIZE-1) & MULT_16_3(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(1,2)(MULT_SIZE-1) & MULT_16_4(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(1,2)<=signed(MULT_16_5(1,2)(MULT_SIZE-1) & MULT_16_5(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(1,2)(MULT_SIZE-1) & MULT_16_6(1,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(1,2) ------------------

			MULTS_1_1_1(1,3)<=signed(MULT_1_1(1,3)(MULT_SIZE-1) & MULT_1_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(1,3)(MULT_SIZE-1) & MULT_1_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(1,3)<=signed(MULT_1_3(1,3)(MULT_SIZE-1) & MULT_1_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(1,3)(MULT_SIZE-1) & MULT_1_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(1,3)<=signed(MULT_1_5(1,3)(MULT_SIZE-1) & MULT_1_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(1,3)(MULT_SIZE-1) & MULT_1_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(1,3)<=signed(MULT_2_1(1,3)(MULT_SIZE-1) & MULT_2_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(1,3)(MULT_SIZE-1) & MULT_2_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(1,3)<=signed(MULT_2_3(1,3)(MULT_SIZE-1) & MULT_2_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(1,3)(MULT_SIZE-1) & MULT_2_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(1,3)<=signed(MULT_2_5(1,3)(MULT_SIZE-1) & MULT_2_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(1,3)(MULT_SIZE-1) & MULT_2_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(1,3)<=signed(MULT_3_1(1,3)(MULT_SIZE-1) & MULT_3_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(1,3)(MULT_SIZE-1) & MULT_3_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(1,3)<=signed(MULT_3_3(1,3)(MULT_SIZE-1) & MULT_3_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(1,3)(MULT_SIZE-1) & MULT_3_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(1,3)<=signed(MULT_3_5(1,3)(MULT_SIZE-1) & MULT_3_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(1,3)(MULT_SIZE-1) & MULT_3_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(1,3)<=signed(MULT_4_1(1,3)(MULT_SIZE-1) & MULT_4_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(1,3)(MULT_SIZE-1) & MULT_4_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(1,3)<=signed(MULT_4_3(1,3)(MULT_SIZE-1) & MULT_4_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(1,3)(MULT_SIZE-1) & MULT_4_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(1,3)<=signed(MULT_4_5(1,3)(MULT_SIZE-1) & MULT_4_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(1,3)(MULT_SIZE-1) & MULT_4_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(1,3)<=signed(MULT_5_1(1,3)(MULT_SIZE-1) & MULT_5_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(1,3)(MULT_SIZE-1) & MULT_5_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(1,3)<=signed(MULT_5_3(1,3)(MULT_SIZE-1) & MULT_5_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(1,3)(MULT_SIZE-1) & MULT_5_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(1,3)<=signed(MULT_5_5(1,3)(MULT_SIZE-1) & MULT_5_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(1,3)(MULT_SIZE-1) & MULT_5_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(1,3)<=signed(MULT_6_1(1,3)(MULT_SIZE-1) & MULT_6_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(1,3)(MULT_SIZE-1) & MULT_6_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(1,3)<=signed(MULT_6_3(1,3)(MULT_SIZE-1) & MULT_6_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(1,3)(MULT_SIZE-1) & MULT_6_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(1,3)<=signed(MULT_6_5(1,3)(MULT_SIZE-1) & MULT_6_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(1,3)(MULT_SIZE-1) & MULT_6_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(1,3)<=signed(MULT_7_1(1,3)(MULT_SIZE-1) & MULT_7_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(1,3)(MULT_SIZE-1) & MULT_7_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(1,3)<=signed(MULT_7_3(1,3)(MULT_SIZE-1) & MULT_7_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(1,3)(MULT_SIZE-1) & MULT_7_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(1,3)<=signed(MULT_7_5(1,3)(MULT_SIZE-1) & MULT_7_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(1,3)(MULT_SIZE-1) & MULT_7_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(1,3)<=signed(MULT_8_1(1,3)(MULT_SIZE-1) & MULT_8_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(1,3)(MULT_SIZE-1) & MULT_8_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(1,3)<=signed(MULT_8_3(1,3)(MULT_SIZE-1) & MULT_8_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(1,3)(MULT_SIZE-1) & MULT_8_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(1,3)<=signed(MULT_8_5(1,3)(MULT_SIZE-1) & MULT_8_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(1,3)(MULT_SIZE-1) & MULT_8_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(1,3)<=signed(MULT_9_1(1,3)(MULT_SIZE-1) & MULT_9_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(1,3)(MULT_SIZE-1) & MULT_9_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(1,3)<=signed(MULT_9_3(1,3)(MULT_SIZE-1) & MULT_9_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(1,3)(MULT_SIZE-1) & MULT_9_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(1,3)<=signed(MULT_9_5(1,3)(MULT_SIZE-1) & MULT_9_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(1,3)(MULT_SIZE-1) & MULT_9_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(1,3)<=signed(MULT_10_1(1,3)(MULT_SIZE-1) & MULT_10_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(1,3)(MULT_SIZE-1) & MULT_10_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(1,3)<=signed(MULT_10_3(1,3)(MULT_SIZE-1) & MULT_10_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(1,3)(MULT_SIZE-1) & MULT_10_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(1,3)<=signed(MULT_10_5(1,3)(MULT_SIZE-1) & MULT_10_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(1,3)(MULT_SIZE-1) & MULT_10_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(1,3)<=signed(MULT_11_1(1,3)(MULT_SIZE-1) & MULT_11_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(1,3)(MULT_SIZE-1) & MULT_11_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(1,3)<=signed(MULT_11_3(1,3)(MULT_SIZE-1) & MULT_11_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(1,3)(MULT_SIZE-1) & MULT_11_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(1,3)<=signed(MULT_11_5(1,3)(MULT_SIZE-1) & MULT_11_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(1,3)(MULT_SIZE-1) & MULT_11_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(1,3)<=signed(MULT_12_1(1,3)(MULT_SIZE-1) & MULT_12_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(1,3)(MULT_SIZE-1) & MULT_12_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(1,3)<=signed(MULT_12_3(1,3)(MULT_SIZE-1) & MULT_12_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(1,3)(MULT_SIZE-1) & MULT_12_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(1,3)<=signed(MULT_12_5(1,3)(MULT_SIZE-1) & MULT_12_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(1,3)(MULT_SIZE-1) & MULT_12_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(1,3)<=signed(MULT_13_1(1,3)(MULT_SIZE-1) & MULT_13_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(1,3)(MULT_SIZE-1) & MULT_13_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(1,3)<=signed(MULT_13_3(1,3)(MULT_SIZE-1) & MULT_13_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(1,3)(MULT_SIZE-1) & MULT_13_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(1,3)<=signed(MULT_13_5(1,3)(MULT_SIZE-1) & MULT_13_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(1,3)(MULT_SIZE-1) & MULT_13_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(1,3)<=signed(MULT_14_1(1,3)(MULT_SIZE-1) & MULT_14_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(1,3)(MULT_SIZE-1) & MULT_14_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(1,3)<=signed(MULT_14_3(1,3)(MULT_SIZE-1) & MULT_14_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(1,3)(MULT_SIZE-1) & MULT_14_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(1,3)<=signed(MULT_14_5(1,3)(MULT_SIZE-1) & MULT_14_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(1,3)(MULT_SIZE-1) & MULT_14_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(1,3)<=signed(MULT_15_1(1,3)(MULT_SIZE-1) & MULT_15_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(1,3)(MULT_SIZE-1) & MULT_15_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(1,3)<=signed(MULT_15_3(1,3)(MULT_SIZE-1) & MULT_15_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(1,3)(MULT_SIZE-1) & MULT_15_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(1,3)<=signed(MULT_15_5(1,3)(MULT_SIZE-1) & MULT_15_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(1,3)(MULT_SIZE-1) & MULT_15_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(1,3)<=signed(MULT_16_1(1,3)(MULT_SIZE-1) & MULT_16_1(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(1,3)(MULT_SIZE-1) & MULT_16_2(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(1,3)<=signed(MULT_16_3(1,3)(MULT_SIZE-1) & MULT_16_3(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(1,3)(MULT_SIZE-1) & MULT_16_4(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(1,3)<=signed(MULT_16_5(1,3)(MULT_SIZE-1) & MULT_16_5(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(1,3)(MULT_SIZE-1) & MULT_16_6(1,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(1,3) ------------------

			MULTS_1_1_1(1,4)<=signed(MULT_1_1(1,4)(MULT_SIZE-1) & MULT_1_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(1,4)(MULT_SIZE-1) & MULT_1_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(1,4)<=signed(MULT_1_3(1,4)(MULT_SIZE-1) & MULT_1_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(1,4)(MULT_SIZE-1) & MULT_1_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(1,4)<=signed(MULT_1_5(1,4)(MULT_SIZE-1) & MULT_1_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(1,4)(MULT_SIZE-1) & MULT_1_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(1,4)<=signed(MULT_2_1(1,4)(MULT_SIZE-1) & MULT_2_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(1,4)(MULT_SIZE-1) & MULT_2_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(1,4)<=signed(MULT_2_3(1,4)(MULT_SIZE-1) & MULT_2_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(1,4)(MULT_SIZE-1) & MULT_2_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(1,4)<=signed(MULT_2_5(1,4)(MULT_SIZE-1) & MULT_2_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(1,4)(MULT_SIZE-1) & MULT_2_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(1,4)<=signed(MULT_3_1(1,4)(MULT_SIZE-1) & MULT_3_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(1,4)(MULT_SIZE-1) & MULT_3_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(1,4)<=signed(MULT_3_3(1,4)(MULT_SIZE-1) & MULT_3_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(1,4)(MULT_SIZE-1) & MULT_3_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(1,4)<=signed(MULT_3_5(1,4)(MULT_SIZE-1) & MULT_3_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(1,4)(MULT_SIZE-1) & MULT_3_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(1,4)<=signed(MULT_4_1(1,4)(MULT_SIZE-1) & MULT_4_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(1,4)(MULT_SIZE-1) & MULT_4_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(1,4)<=signed(MULT_4_3(1,4)(MULT_SIZE-1) & MULT_4_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(1,4)(MULT_SIZE-1) & MULT_4_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(1,4)<=signed(MULT_4_5(1,4)(MULT_SIZE-1) & MULT_4_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(1,4)(MULT_SIZE-1) & MULT_4_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(1,4)<=signed(MULT_5_1(1,4)(MULT_SIZE-1) & MULT_5_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(1,4)(MULT_SIZE-1) & MULT_5_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(1,4)<=signed(MULT_5_3(1,4)(MULT_SIZE-1) & MULT_5_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(1,4)(MULT_SIZE-1) & MULT_5_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(1,4)<=signed(MULT_5_5(1,4)(MULT_SIZE-1) & MULT_5_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(1,4)(MULT_SIZE-1) & MULT_5_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(1,4)<=signed(MULT_6_1(1,4)(MULT_SIZE-1) & MULT_6_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(1,4)(MULT_SIZE-1) & MULT_6_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(1,4)<=signed(MULT_6_3(1,4)(MULT_SIZE-1) & MULT_6_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(1,4)(MULT_SIZE-1) & MULT_6_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(1,4)<=signed(MULT_6_5(1,4)(MULT_SIZE-1) & MULT_6_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(1,4)(MULT_SIZE-1) & MULT_6_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(1,4)<=signed(MULT_7_1(1,4)(MULT_SIZE-1) & MULT_7_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(1,4)(MULT_SIZE-1) & MULT_7_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(1,4)<=signed(MULT_7_3(1,4)(MULT_SIZE-1) & MULT_7_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(1,4)(MULT_SIZE-1) & MULT_7_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(1,4)<=signed(MULT_7_5(1,4)(MULT_SIZE-1) & MULT_7_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(1,4)(MULT_SIZE-1) & MULT_7_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(1,4)<=signed(MULT_8_1(1,4)(MULT_SIZE-1) & MULT_8_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(1,4)(MULT_SIZE-1) & MULT_8_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(1,4)<=signed(MULT_8_3(1,4)(MULT_SIZE-1) & MULT_8_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(1,4)(MULT_SIZE-1) & MULT_8_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(1,4)<=signed(MULT_8_5(1,4)(MULT_SIZE-1) & MULT_8_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(1,4)(MULT_SIZE-1) & MULT_8_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(1,4)<=signed(MULT_9_1(1,4)(MULT_SIZE-1) & MULT_9_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(1,4)(MULT_SIZE-1) & MULT_9_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(1,4)<=signed(MULT_9_3(1,4)(MULT_SIZE-1) & MULT_9_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(1,4)(MULT_SIZE-1) & MULT_9_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(1,4)<=signed(MULT_9_5(1,4)(MULT_SIZE-1) & MULT_9_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(1,4)(MULT_SIZE-1) & MULT_9_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(1,4)<=signed(MULT_10_1(1,4)(MULT_SIZE-1) & MULT_10_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(1,4)(MULT_SIZE-1) & MULT_10_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(1,4)<=signed(MULT_10_3(1,4)(MULT_SIZE-1) & MULT_10_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(1,4)(MULT_SIZE-1) & MULT_10_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(1,4)<=signed(MULT_10_5(1,4)(MULT_SIZE-1) & MULT_10_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(1,4)(MULT_SIZE-1) & MULT_10_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(1,4)<=signed(MULT_11_1(1,4)(MULT_SIZE-1) & MULT_11_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(1,4)(MULT_SIZE-1) & MULT_11_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(1,4)<=signed(MULT_11_3(1,4)(MULT_SIZE-1) & MULT_11_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(1,4)(MULT_SIZE-1) & MULT_11_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(1,4)<=signed(MULT_11_5(1,4)(MULT_SIZE-1) & MULT_11_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(1,4)(MULT_SIZE-1) & MULT_11_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(1,4)<=signed(MULT_12_1(1,4)(MULT_SIZE-1) & MULT_12_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(1,4)(MULT_SIZE-1) & MULT_12_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(1,4)<=signed(MULT_12_3(1,4)(MULT_SIZE-1) & MULT_12_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(1,4)(MULT_SIZE-1) & MULT_12_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(1,4)<=signed(MULT_12_5(1,4)(MULT_SIZE-1) & MULT_12_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(1,4)(MULT_SIZE-1) & MULT_12_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(1,4)<=signed(MULT_13_1(1,4)(MULT_SIZE-1) & MULT_13_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(1,4)(MULT_SIZE-1) & MULT_13_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(1,4)<=signed(MULT_13_3(1,4)(MULT_SIZE-1) & MULT_13_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(1,4)(MULT_SIZE-1) & MULT_13_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(1,4)<=signed(MULT_13_5(1,4)(MULT_SIZE-1) & MULT_13_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(1,4)(MULT_SIZE-1) & MULT_13_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(1,4)<=signed(MULT_14_1(1,4)(MULT_SIZE-1) & MULT_14_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(1,4)(MULT_SIZE-1) & MULT_14_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(1,4)<=signed(MULT_14_3(1,4)(MULT_SIZE-1) & MULT_14_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(1,4)(MULT_SIZE-1) & MULT_14_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(1,4)<=signed(MULT_14_5(1,4)(MULT_SIZE-1) & MULT_14_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(1,4)(MULT_SIZE-1) & MULT_14_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(1,4)<=signed(MULT_15_1(1,4)(MULT_SIZE-1) & MULT_15_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(1,4)(MULT_SIZE-1) & MULT_15_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(1,4)<=signed(MULT_15_3(1,4)(MULT_SIZE-1) & MULT_15_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(1,4)(MULT_SIZE-1) & MULT_15_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(1,4)<=signed(MULT_15_5(1,4)(MULT_SIZE-1) & MULT_15_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(1,4)(MULT_SIZE-1) & MULT_15_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(1,4)<=signed(MULT_16_1(1,4)(MULT_SIZE-1) & MULT_16_1(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(1,4)(MULT_SIZE-1) & MULT_16_2(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(1,4)<=signed(MULT_16_3(1,4)(MULT_SIZE-1) & MULT_16_3(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(1,4)(MULT_SIZE-1) & MULT_16_4(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(1,4)<=signed(MULT_16_5(1,4)(MULT_SIZE-1) & MULT_16_5(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(1,4)(MULT_SIZE-1) & MULT_16_6(1,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(1,4) ------------------

			MULTS_1_1_1(2,0)<=signed(MULT_1_1(2,0)(MULT_SIZE-1) & MULT_1_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(2,0)(MULT_SIZE-1) & MULT_1_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(2,0)<=signed(MULT_1_3(2,0)(MULT_SIZE-1) & MULT_1_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(2,0)(MULT_SIZE-1) & MULT_1_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(2,0)<=signed(MULT_1_5(2,0)(MULT_SIZE-1) & MULT_1_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(2,0)(MULT_SIZE-1) & MULT_1_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(2,0)<=signed(MULT_2_1(2,0)(MULT_SIZE-1) & MULT_2_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(2,0)(MULT_SIZE-1) & MULT_2_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(2,0)<=signed(MULT_2_3(2,0)(MULT_SIZE-1) & MULT_2_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(2,0)(MULT_SIZE-1) & MULT_2_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(2,0)<=signed(MULT_2_5(2,0)(MULT_SIZE-1) & MULT_2_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(2,0)(MULT_SIZE-1) & MULT_2_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(2,0)<=signed(MULT_3_1(2,0)(MULT_SIZE-1) & MULT_3_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(2,0)(MULT_SIZE-1) & MULT_3_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(2,0)<=signed(MULT_3_3(2,0)(MULT_SIZE-1) & MULT_3_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(2,0)(MULT_SIZE-1) & MULT_3_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(2,0)<=signed(MULT_3_5(2,0)(MULT_SIZE-1) & MULT_3_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(2,0)(MULT_SIZE-1) & MULT_3_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(2,0)<=signed(MULT_4_1(2,0)(MULT_SIZE-1) & MULT_4_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(2,0)(MULT_SIZE-1) & MULT_4_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(2,0)<=signed(MULT_4_3(2,0)(MULT_SIZE-1) & MULT_4_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(2,0)(MULT_SIZE-1) & MULT_4_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(2,0)<=signed(MULT_4_5(2,0)(MULT_SIZE-1) & MULT_4_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(2,0)(MULT_SIZE-1) & MULT_4_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(2,0)<=signed(MULT_5_1(2,0)(MULT_SIZE-1) & MULT_5_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(2,0)(MULT_SIZE-1) & MULT_5_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(2,0)<=signed(MULT_5_3(2,0)(MULT_SIZE-1) & MULT_5_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(2,0)(MULT_SIZE-1) & MULT_5_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(2,0)<=signed(MULT_5_5(2,0)(MULT_SIZE-1) & MULT_5_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(2,0)(MULT_SIZE-1) & MULT_5_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(2,0)<=signed(MULT_6_1(2,0)(MULT_SIZE-1) & MULT_6_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(2,0)(MULT_SIZE-1) & MULT_6_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(2,0)<=signed(MULT_6_3(2,0)(MULT_SIZE-1) & MULT_6_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(2,0)(MULT_SIZE-1) & MULT_6_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(2,0)<=signed(MULT_6_5(2,0)(MULT_SIZE-1) & MULT_6_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(2,0)(MULT_SIZE-1) & MULT_6_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(2,0)<=signed(MULT_7_1(2,0)(MULT_SIZE-1) & MULT_7_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(2,0)(MULT_SIZE-1) & MULT_7_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(2,0)<=signed(MULT_7_3(2,0)(MULT_SIZE-1) & MULT_7_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(2,0)(MULT_SIZE-1) & MULT_7_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(2,0)<=signed(MULT_7_5(2,0)(MULT_SIZE-1) & MULT_7_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(2,0)(MULT_SIZE-1) & MULT_7_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(2,0)<=signed(MULT_8_1(2,0)(MULT_SIZE-1) & MULT_8_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(2,0)(MULT_SIZE-1) & MULT_8_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(2,0)<=signed(MULT_8_3(2,0)(MULT_SIZE-1) & MULT_8_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(2,0)(MULT_SIZE-1) & MULT_8_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(2,0)<=signed(MULT_8_5(2,0)(MULT_SIZE-1) & MULT_8_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(2,0)(MULT_SIZE-1) & MULT_8_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(2,0)<=signed(MULT_9_1(2,0)(MULT_SIZE-1) & MULT_9_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(2,0)(MULT_SIZE-1) & MULT_9_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(2,0)<=signed(MULT_9_3(2,0)(MULT_SIZE-1) & MULT_9_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(2,0)(MULT_SIZE-1) & MULT_9_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(2,0)<=signed(MULT_9_5(2,0)(MULT_SIZE-1) & MULT_9_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(2,0)(MULT_SIZE-1) & MULT_9_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(2,0)<=signed(MULT_10_1(2,0)(MULT_SIZE-1) & MULT_10_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(2,0)(MULT_SIZE-1) & MULT_10_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(2,0)<=signed(MULT_10_3(2,0)(MULT_SIZE-1) & MULT_10_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(2,0)(MULT_SIZE-1) & MULT_10_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(2,0)<=signed(MULT_10_5(2,0)(MULT_SIZE-1) & MULT_10_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(2,0)(MULT_SIZE-1) & MULT_10_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(2,0)<=signed(MULT_11_1(2,0)(MULT_SIZE-1) & MULT_11_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(2,0)(MULT_SIZE-1) & MULT_11_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(2,0)<=signed(MULT_11_3(2,0)(MULT_SIZE-1) & MULT_11_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(2,0)(MULT_SIZE-1) & MULT_11_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(2,0)<=signed(MULT_11_5(2,0)(MULT_SIZE-1) & MULT_11_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(2,0)(MULT_SIZE-1) & MULT_11_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(2,0)<=signed(MULT_12_1(2,0)(MULT_SIZE-1) & MULT_12_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(2,0)(MULT_SIZE-1) & MULT_12_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(2,0)<=signed(MULT_12_3(2,0)(MULT_SIZE-1) & MULT_12_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(2,0)(MULT_SIZE-1) & MULT_12_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(2,0)<=signed(MULT_12_5(2,0)(MULT_SIZE-1) & MULT_12_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(2,0)(MULT_SIZE-1) & MULT_12_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(2,0)<=signed(MULT_13_1(2,0)(MULT_SIZE-1) & MULT_13_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(2,0)(MULT_SIZE-1) & MULT_13_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(2,0)<=signed(MULT_13_3(2,0)(MULT_SIZE-1) & MULT_13_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(2,0)(MULT_SIZE-1) & MULT_13_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(2,0)<=signed(MULT_13_5(2,0)(MULT_SIZE-1) & MULT_13_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(2,0)(MULT_SIZE-1) & MULT_13_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(2,0)<=signed(MULT_14_1(2,0)(MULT_SIZE-1) & MULT_14_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(2,0)(MULT_SIZE-1) & MULT_14_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(2,0)<=signed(MULT_14_3(2,0)(MULT_SIZE-1) & MULT_14_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(2,0)(MULT_SIZE-1) & MULT_14_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(2,0)<=signed(MULT_14_5(2,0)(MULT_SIZE-1) & MULT_14_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(2,0)(MULT_SIZE-1) & MULT_14_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(2,0)<=signed(MULT_15_1(2,0)(MULT_SIZE-1) & MULT_15_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(2,0)(MULT_SIZE-1) & MULT_15_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(2,0)<=signed(MULT_15_3(2,0)(MULT_SIZE-1) & MULT_15_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(2,0)(MULT_SIZE-1) & MULT_15_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(2,0)<=signed(MULT_15_5(2,0)(MULT_SIZE-1) & MULT_15_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(2,0)(MULT_SIZE-1) & MULT_15_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(2,0)<=signed(MULT_16_1(2,0)(MULT_SIZE-1) & MULT_16_1(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(2,0)(MULT_SIZE-1) & MULT_16_2(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(2,0)<=signed(MULT_16_3(2,0)(MULT_SIZE-1) & MULT_16_3(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(2,0)(MULT_SIZE-1) & MULT_16_4(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(2,0)<=signed(MULT_16_5(2,0)(MULT_SIZE-1) & MULT_16_5(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(2,0)(MULT_SIZE-1) & MULT_16_6(2,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(2,0) ------------------

			MULTS_1_1_1(2,1)<=signed(MULT_1_1(2,1)(MULT_SIZE-1) & MULT_1_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(2,1)(MULT_SIZE-1) & MULT_1_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(2,1)<=signed(MULT_1_3(2,1)(MULT_SIZE-1) & MULT_1_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(2,1)(MULT_SIZE-1) & MULT_1_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(2,1)<=signed(MULT_1_5(2,1)(MULT_SIZE-1) & MULT_1_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(2,1)(MULT_SIZE-1) & MULT_1_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(2,1)<=signed(MULT_2_1(2,1)(MULT_SIZE-1) & MULT_2_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(2,1)(MULT_SIZE-1) & MULT_2_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(2,1)<=signed(MULT_2_3(2,1)(MULT_SIZE-1) & MULT_2_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(2,1)(MULT_SIZE-1) & MULT_2_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(2,1)<=signed(MULT_2_5(2,1)(MULT_SIZE-1) & MULT_2_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(2,1)(MULT_SIZE-1) & MULT_2_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(2,1)<=signed(MULT_3_1(2,1)(MULT_SIZE-1) & MULT_3_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(2,1)(MULT_SIZE-1) & MULT_3_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(2,1)<=signed(MULT_3_3(2,1)(MULT_SIZE-1) & MULT_3_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(2,1)(MULT_SIZE-1) & MULT_3_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(2,1)<=signed(MULT_3_5(2,1)(MULT_SIZE-1) & MULT_3_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(2,1)(MULT_SIZE-1) & MULT_3_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(2,1)<=signed(MULT_4_1(2,1)(MULT_SIZE-1) & MULT_4_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(2,1)(MULT_SIZE-1) & MULT_4_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(2,1)<=signed(MULT_4_3(2,1)(MULT_SIZE-1) & MULT_4_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(2,1)(MULT_SIZE-1) & MULT_4_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(2,1)<=signed(MULT_4_5(2,1)(MULT_SIZE-1) & MULT_4_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(2,1)(MULT_SIZE-1) & MULT_4_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(2,1)<=signed(MULT_5_1(2,1)(MULT_SIZE-1) & MULT_5_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(2,1)(MULT_SIZE-1) & MULT_5_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(2,1)<=signed(MULT_5_3(2,1)(MULT_SIZE-1) & MULT_5_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(2,1)(MULT_SIZE-1) & MULT_5_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(2,1)<=signed(MULT_5_5(2,1)(MULT_SIZE-1) & MULT_5_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(2,1)(MULT_SIZE-1) & MULT_5_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(2,1)<=signed(MULT_6_1(2,1)(MULT_SIZE-1) & MULT_6_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(2,1)(MULT_SIZE-1) & MULT_6_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(2,1)<=signed(MULT_6_3(2,1)(MULT_SIZE-1) & MULT_6_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(2,1)(MULT_SIZE-1) & MULT_6_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(2,1)<=signed(MULT_6_5(2,1)(MULT_SIZE-1) & MULT_6_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(2,1)(MULT_SIZE-1) & MULT_6_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(2,1)<=signed(MULT_7_1(2,1)(MULT_SIZE-1) & MULT_7_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(2,1)(MULT_SIZE-1) & MULT_7_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(2,1)<=signed(MULT_7_3(2,1)(MULT_SIZE-1) & MULT_7_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(2,1)(MULT_SIZE-1) & MULT_7_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(2,1)<=signed(MULT_7_5(2,1)(MULT_SIZE-1) & MULT_7_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(2,1)(MULT_SIZE-1) & MULT_7_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(2,1)<=signed(MULT_8_1(2,1)(MULT_SIZE-1) & MULT_8_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(2,1)(MULT_SIZE-1) & MULT_8_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(2,1)<=signed(MULT_8_3(2,1)(MULT_SIZE-1) & MULT_8_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(2,1)(MULT_SIZE-1) & MULT_8_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(2,1)<=signed(MULT_8_5(2,1)(MULT_SIZE-1) & MULT_8_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(2,1)(MULT_SIZE-1) & MULT_8_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(2,1)<=signed(MULT_9_1(2,1)(MULT_SIZE-1) & MULT_9_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(2,1)(MULT_SIZE-1) & MULT_9_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(2,1)<=signed(MULT_9_3(2,1)(MULT_SIZE-1) & MULT_9_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(2,1)(MULT_SIZE-1) & MULT_9_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(2,1)<=signed(MULT_9_5(2,1)(MULT_SIZE-1) & MULT_9_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(2,1)(MULT_SIZE-1) & MULT_9_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(2,1)<=signed(MULT_10_1(2,1)(MULT_SIZE-1) & MULT_10_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(2,1)(MULT_SIZE-1) & MULT_10_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(2,1)<=signed(MULT_10_3(2,1)(MULT_SIZE-1) & MULT_10_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(2,1)(MULT_SIZE-1) & MULT_10_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(2,1)<=signed(MULT_10_5(2,1)(MULT_SIZE-1) & MULT_10_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(2,1)(MULT_SIZE-1) & MULT_10_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(2,1)<=signed(MULT_11_1(2,1)(MULT_SIZE-1) & MULT_11_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(2,1)(MULT_SIZE-1) & MULT_11_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(2,1)<=signed(MULT_11_3(2,1)(MULT_SIZE-1) & MULT_11_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(2,1)(MULT_SIZE-1) & MULT_11_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(2,1)<=signed(MULT_11_5(2,1)(MULT_SIZE-1) & MULT_11_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(2,1)(MULT_SIZE-1) & MULT_11_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(2,1)<=signed(MULT_12_1(2,1)(MULT_SIZE-1) & MULT_12_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(2,1)(MULT_SIZE-1) & MULT_12_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(2,1)<=signed(MULT_12_3(2,1)(MULT_SIZE-1) & MULT_12_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(2,1)(MULT_SIZE-1) & MULT_12_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(2,1)<=signed(MULT_12_5(2,1)(MULT_SIZE-1) & MULT_12_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(2,1)(MULT_SIZE-1) & MULT_12_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(2,1)<=signed(MULT_13_1(2,1)(MULT_SIZE-1) & MULT_13_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(2,1)(MULT_SIZE-1) & MULT_13_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(2,1)<=signed(MULT_13_3(2,1)(MULT_SIZE-1) & MULT_13_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(2,1)(MULT_SIZE-1) & MULT_13_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(2,1)<=signed(MULT_13_5(2,1)(MULT_SIZE-1) & MULT_13_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(2,1)(MULT_SIZE-1) & MULT_13_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(2,1)<=signed(MULT_14_1(2,1)(MULT_SIZE-1) & MULT_14_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(2,1)(MULT_SIZE-1) & MULT_14_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(2,1)<=signed(MULT_14_3(2,1)(MULT_SIZE-1) & MULT_14_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(2,1)(MULT_SIZE-1) & MULT_14_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(2,1)<=signed(MULT_14_5(2,1)(MULT_SIZE-1) & MULT_14_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(2,1)(MULT_SIZE-1) & MULT_14_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(2,1)<=signed(MULT_15_1(2,1)(MULT_SIZE-1) & MULT_15_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(2,1)(MULT_SIZE-1) & MULT_15_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(2,1)<=signed(MULT_15_3(2,1)(MULT_SIZE-1) & MULT_15_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(2,1)(MULT_SIZE-1) & MULT_15_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(2,1)<=signed(MULT_15_5(2,1)(MULT_SIZE-1) & MULT_15_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(2,1)(MULT_SIZE-1) & MULT_15_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(2,1)<=signed(MULT_16_1(2,1)(MULT_SIZE-1) & MULT_16_1(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(2,1)(MULT_SIZE-1) & MULT_16_2(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(2,1)<=signed(MULT_16_3(2,1)(MULT_SIZE-1) & MULT_16_3(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(2,1)(MULT_SIZE-1) & MULT_16_4(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(2,1)<=signed(MULT_16_5(2,1)(MULT_SIZE-1) & MULT_16_5(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(2,1)(MULT_SIZE-1) & MULT_16_6(2,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(2,1) ------------------

			MULTS_1_1_1(2,2)<=signed(MULT_1_1(2,2)(MULT_SIZE-1) & MULT_1_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(2,2)(MULT_SIZE-1) & MULT_1_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(2,2)<=signed(MULT_1_3(2,2)(MULT_SIZE-1) & MULT_1_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(2,2)(MULT_SIZE-1) & MULT_1_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(2,2)<=signed(MULT_1_5(2,2)(MULT_SIZE-1) & MULT_1_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(2,2)(MULT_SIZE-1) & MULT_1_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(2,2)<=signed(MULT_2_1(2,2)(MULT_SIZE-1) & MULT_2_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(2,2)(MULT_SIZE-1) & MULT_2_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(2,2)<=signed(MULT_2_3(2,2)(MULT_SIZE-1) & MULT_2_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(2,2)(MULT_SIZE-1) & MULT_2_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(2,2)<=signed(MULT_2_5(2,2)(MULT_SIZE-1) & MULT_2_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(2,2)(MULT_SIZE-1) & MULT_2_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(2,2)<=signed(MULT_3_1(2,2)(MULT_SIZE-1) & MULT_3_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(2,2)(MULT_SIZE-1) & MULT_3_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(2,2)<=signed(MULT_3_3(2,2)(MULT_SIZE-1) & MULT_3_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(2,2)(MULT_SIZE-1) & MULT_3_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(2,2)<=signed(MULT_3_5(2,2)(MULT_SIZE-1) & MULT_3_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(2,2)(MULT_SIZE-1) & MULT_3_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(2,2)<=signed(MULT_4_1(2,2)(MULT_SIZE-1) & MULT_4_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(2,2)(MULT_SIZE-1) & MULT_4_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(2,2)<=signed(MULT_4_3(2,2)(MULT_SIZE-1) & MULT_4_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(2,2)(MULT_SIZE-1) & MULT_4_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(2,2)<=signed(MULT_4_5(2,2)(MULT_SIZE-1) & MULT_4_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(2,2)(MULT_SIZE-1) & MULT_4_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(2,2)<=signed(MULT_5_1(2,2)(MULT_SIZE-1) & MULT_5_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(2,2)(MULT_SIZE-1) & MULT_5_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(2,2)<=signed(MULT_5_3(2,2)(MULT_SIZE-1) & MULT_5_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(2,2)(MULT_SIZE-1) & MULT_5_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(2,2)<=signed(MULT_5_5(2,2)(MULT_SIZE-1) & MULT_5_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(2,2)(MULT_SIZE-1) & MULT_5_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(2,2)<=signed(MULT_6_1(2,2)(MULT_SIZE-1) & MULT_6_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(2,2)(MULT_SIZE-1) & MULT_6_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(2,2)<=signed(MULT_6_3(2,2)(MULT_SIZE-1) & MULT_6_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(2,2)(MULT_SIZE-1) & MULT_6_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(2,2)<=signed(MULT_6_5(2,2)(MULT_SIZE-1) & MULT_6_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(2,2)(MULT_SIZE-1) & MULT_6_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(2,2)<=signed(MULT_7_1(2,2)(MULT_SIZE-1) & MULT_7_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(2,2)(MULT_SIZE-1) & MULT_7_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(2,2)<=signed(MULT_7_3(2,2)(MULT_SIZE-1) & MULT_7_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(2,2)(MULT_SIZE-1) & MULT_7_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(2,2)<=signed(MULT_7_5(2,2)(MULT_SIZE-1) & MULT_7_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(2,2)(MULT_SIZE-1) & MULT_7_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(2,2)<=signed(MULT_8_1(2,2)(MULT_SIZE-1) & MULT_8_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(2,2)(MULT_SIZE-1) & MULT_8_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(2,2)<=signed(MULT_8_3(2,2)(MULT_SIZE-1) & MULT_8_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(2,2)(MULT_SIZE-1) & MULT_8_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(2,2)<=signed(MULT_8_5(2,2)(MULT_SIZE-1) & MULT_8_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(2,2)(MULT_SIZE-1) & MULT_8_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(2,2)<=signed(MULT_9_1(2,2)(MULT_SIZE-1) & MULT_9_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(2,2)(MULT_SIZE-1) & MULT_9_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(2,2)<=signed(MULT_9_3(2,2)(MULT_SIZE-1) & MULT_9_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(2,2)(MULT_SIZE-1) & MULT_9_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(2,2)<=signed(MULT_9_5(2,2)(MULT_SIZE-1) & MULT_9_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(2,2)(MULT_SIZE-1) & MULT_9_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(2,2)<=signed(MULT_10_1(2,2)(MULT_SIZE-1) & MULT_10_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(2,2)(MULT_SIZE-1) & MULT_10_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(2,2)<=signed(MULT_10_3(2,2)(MULT_SIZE-1) & MULT_10_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(2,2)(MULT_SIZE-1) & MULT_10_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(2,2)<=signed(MULT_10_5(2,2)(MULT_SIZE-1) & MULT_10_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(2,2)(MULT_SIZE-1) & MULT_10_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(2,2)<=signed(MULT_11_1(2,2)(MULT_SIZE-1) & MULT_11_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(2,2)(MULT_SIZE-1) & MULT_11_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(2,2)<=signed(MULT_11_3(2,2)(MULT_SIZE-1) & MULT_11_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(2,2)(MULT_SIZE-1) & MULT_11_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(2,2)<=signed(MULT_11_5(2,2)(MULT_SIZE-1) & MULT_11_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(2,2)(MULT_SIZE-1) & MULT_11_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(2,2)<=signed(MULT_12_1(2,2)(MULT_SIZE-1) & MULT_12_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(2,2)(MULT_SIZE-1) & MULT_12_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(2,2)<=signed(MULT_12_3(2,2)(MULT_SIZE-1) & MULT_12_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(2,2)(MULT_SIZE-1) & MULT_12_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(2,2)<=signed(MULT_12_5(2,2)(MULT_SIZE-1) & MULT_12_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(2,2)(MULT_SIZE-1) & MULT_12_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(2,2)<=signed(MULT_13_1(2,2)(MULT_SIZE-1) & MULT_13_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(2,2)(MULT_SIZE-1) & MULT_13_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(2,2)<=signed(MULT_13_3(2,2)(MULT_SIZE-1) & MULT_13_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(2,2)(MULT_SIZE-1) & MULT_13_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(2,2)<=signed(MULT_13_5(2,2)(MULT_SIZE-1) & MULT_13_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(2,2)(MULT_SIZE-1) & MULT_13_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(2,2)<=signed(MULT_14_1(2,2)(MULT_SIZE-1) & MULT_14_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(2,2)(MULT_SIZE-1) & MULT_14_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(2,2)<=signed(MULT_14_3(2,2)(MULT_SIZE-1) & MULT_14_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(2,2)(MULT_SIZE-1) & MULT_14_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(2,2)<=signed(MULT_14_5(2,2)(MULT_SIZE-1) & MULT_14_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(2,2)(MULT_SIZE-1) & MULT_14_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(2,2)<=signed(MULT_15_1(2,2)(MULT_SIZE-1) & MULT_15_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(2,2)(MULT_SIZE-1) & MULT_15_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(2,2)<=signed(MULT_15_3(2,2)(MULT_SIZE-1) & MULT_15_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(2,2)(MULT_SIZE-1) & MULT_15_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(2,2)<=signed(MULT_15_5(2,2)(MULT_SIZE-1) & MULT_15_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(2,2)(MULT_SIZE-1) & MULT_15_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(2,2)<=signed(MULT_16_1(2,2)(MULT_SIZE-1) & MULT_16_1(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(2,2)(MULT_SIZE-1) & MULT_16_2(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(2,2)<=signed(MULT_16_3(2,2)(MULT_SIZE-1) & MULT_16_3(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(2,2)(MULT_SIZE-1) & MULT_16_4(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(2,2)<=signed(MULT_16_5(2,2)(MULT_SIZE-1) & MULT_16_5(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(2,2)(MULT_SIZE-1) & MULT_16_6(2,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(2,2) ------------------

			MULTS_1_1_1(2,3)<=signed(MULT_1_1(2,3)(MULT_SIZE-1) & MULT_1_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(2,3)(MULT_SIZE-1) & MULT_1_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(2,3)<=signed(MULT_1_3(2,3)(MULT_SIZE-1) & MULT_1_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(2,3)(MULT_SIZE-1) & MULT_1_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(2,3)<=signed(MULT_1_5(2,3)(MULT_SIZE-1) & MULT_1_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(2,3)(MULT_SIZE-1) & MULT_1_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(2,3)<=signed(MULT_2_1(2,3)(MULT_SIZE-1) & MULT_2_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(2,3)(MULT_SIZE-1) & MULT_2_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(2,3)<=signed(MULT_2_3(2,3)(MULT_SIZE-1) & MULT_2_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(2,3)(MULT_SIZE-1) & MULT_2_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(2,3)<=signed(MULT_2_5(2,3)(MULT_SIZE-1) & MULT_2_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(2,3)(MULT_SIZE-1) & MULT_2_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(2,3)<=signed(MULT_3_1(2,3)(MULT_SIZE-1) & MULT_3_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(2,3)(MULT_SIZE-1) & MULT_3_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(2,3)<=signed(MULT_3_3(2,3)(MULT_SIZE-1) & MULT_3_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(2,3)(MULT_SIZE-1) & MULT_3_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(2,3)<=signed(MULT_3_5(2,3)(MULT_SIZE-1) & MULT_3_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(2,3)(MULT_SIZE-1) & MULT_3_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(2,3)<=signed(MULT_4_1(2,3)(MULT_SIZE-1) & MULT_4_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(2,3)(MULT_SIZE-1) & MULT_4_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(2,3)<=signed(MULT_4_3(2,3)(MULT_SIZE-1) & MULT_4_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(2,3)(MULT_SIZE-1) & MULT_4_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(2,3)<=signed(MULT_4_5(2,3)(MULT_SIZE-1) & MULT_4_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(2,3)(MULT_SIZE-1) & MULT_4_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(2,3)<=signed(MULT_5_1(2,3)(MULT_SIZE-1) & MULT_5_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(2,3)(MULT_SIZE-1) & MULT_5_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(2,3)<=signed(MULT_5_3(2,3)(MULT_SIZE-1) & MULT_5_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(2,3)(MULT_SIZE-1) & MULT_5_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(2,3)<=signed(MULT_5_5(2,3)(MULT_SIZE-1) & MULT_5_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(2,3)(MULT_SIZE-1) & MULT_5_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(2,3)<=signed(MULT_6_1(2,3)(MULT_SIZE-1) & MULT_6_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(2,3)(MULT_SIZE-1) & MULT_6_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(2,3)<=signed(MULT_6_3(2,3)(MULT_SIZE-1) & MULT_6_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(2,3)(MULT_SIZE-1) & MULT_6_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(2,3)<=signed(MULT_6_5(2,3)(MULT_SIZE-1) & MULT_6_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(2,3)(MULT_SIZE-1) & MULT_6_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(2,3)<=signed(MULT_7_1(2,3)(MULT_SIZE-1) & MULT_7_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(2,3)(MULT_SIZE-1) & MULT_7_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(2,3)<=signed(MULT_7_3(2,3)(MULT_SIZE-1) & MULT_7_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(2,3)(MULT_SIZE-1) & MULT_7_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(2,3)<=signed(MULT_7_5(2,3)(MULT_SIZE-1) & MULT_7_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(2,3)(MULT_SIZE-1) & MULT_7_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(2,3)<=signed(MULT_8_1(2,3)(MULT_SIZE-1) & MULT_8_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(2,3)(MULT_SIZE-1) & MULT_8_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(2,3)<=signed(MULT_8_3(2,3)(MULT_SIZE-1) & MULT_8_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(2,3)(MULT_SIZE-1) & MULT_8_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(2,3)<=signed(MULT_8_5(2,3)(MULT_SIZE-1) & MULT_8_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(2,3)(MULT_SIZE-1) & MULT_8_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(2,3)<=signed(MULT_9_1(2,3)(MULT_SIZE-1) & MULT_9_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(2,3)(MULT_SIZE-1) & MULT_9_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(2,3)<=signed(MULT_9_3(2,3)(MULT_SIZE-1) & MULT_9_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(2,3)(MULT_SIZE-1) & MULT_9_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(2,3)<=signed(MULT_9_5(2,3)(MULT_SIZE-1) & MULT_9_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(2,3)(MULT_SIZE-1) & MULT_9_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(2,3)<=signed(MULT_10_1(2,3)(MULT_SIZE-1) & MULT_10_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(2,3)(MULT_SIZE-1) & MULT_10_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(2,3)<=signed(MULT_10_3(2,3)(MULT_SIZE-1) & MULT_10_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(2,3)(MULT_SIZE-1) & MULT_10_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(2,3)<=signed(MULT_10_5(2,3)(MULT_SIZE-1) & MULT_10_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(2,3)(MULT_SIZE-1) & MULT_10_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(2,3)<=signed(MULT_11_1(2,3)(MULT_SIZE-1) & MULT_11_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(2,3)(MULT_SIZE-1) & MULT_11_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(2,3)<=signed(MULT_11_3(2,3)(MULT_SIZE-1) & MULT_11_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(2,3)(MULT_SIZE-1) & MULT_11_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(2,3)<=signed(MULT_11_5(2,3)(MULT_SIZE-1) & MULT_11_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(2,3)(MULT_SIZE-1) & MULT_11_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(2,3)<=signed(MULT_12_1(2,3)(MULT_SIZE-1) & MULT_12_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(2,3)(MULT_SIZE-1) & MULT_12_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(2,3)<=signed(MULT_12_3(2,3)(MULT_SIZE-1) & MULT_12_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(2,3)(MULT_SIZE-1) & MULT_12_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(2,3)<=signed(MULT_12_5(2,3)(MULT_SIZE-1) & MULT_12_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(2,3)(MULT_SIZE-1) & MULT_12_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(2,3)<=signed(MULT_13_1(2,3)(MULT_SIZE-1) & MULT_13_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(2,3)(MULT_SIZE-1) & MULT_13_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(2,3)<=signed(MULT_13_3(2,3)(MULT_SIZE-1) & MULT_13_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(2,3)(MULT_SIZE-1) & MULT_13_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(2,3)<=signed(MULT_13_5(2,3)(MULT_SIZE-1) & MULT_13_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(2,3)(MULT_SIZE-1) & MULT_13_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(2,3)<=signed(MULT_14_1(2,3)(MULT_SIZE-1) & MULT_14_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(2,3)(MULT_SIZE-1) & MULT_14_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(2,3)<=signed(MULT_14_3(2,3)(MULT_SIZE-1) & MULT_14_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(2,3)(MULT_SIZE-1) & MULT_14_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(2,3)<=signed(MULT_14_5(2,3)(MULT_SIZE-1) & MULT_14_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(2,3)(MULT_SIZE-1) & MULT_14_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(2,3)<=signed(MULT_15_1(2,3)(MULT_SIZE-1) & MULT_15_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(2,3)(MULT_SIZE-1) & MULT_15_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(2,3)<=signed(MULT_15_3(2,3)(MULT_SIZE-1) & MULT_15_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(2,3)(MULT_SIZE-1) & MULT_15_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(2,3)<=signed(MULT_15_5(2,3)(MULT_SIZE-1) & MULT_15_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(2,3)(MULT_SIZE-1) & MULT_15_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(2,3)<=signed(MULT_16_1(2,3)(MULT_SIZE-1) & MULT_16_1(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(2,3)(MULT_SIZE-1) & MULT_16_2(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(2,3)<=signed(MULT_16_3(2,3)(MULT_SIZE-1) & MULT_16_3(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(2,3)(MULT_SIZE-1) & MULT_16_4(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(2,3)<=signed(MULT_16_5(2,3)(MULT_SIZE-1) & MULT_16_5(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(2,3)(MULT_SIZE-1) & MULT_16_6(2,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(2,3) ------------------

			MULTS_1_1_1(2,4)<=signed(MULT_1_1(2,4)(MULT_SIZE-1) & MULT_1_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(2,4)(MULT_SIZE-1) & MULT_1_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(2,4)<=signed(MULT_1_3(2,4)(MULT_SIZE-1) & MULT_1_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(2,4)(MULT_SIZE-1) & MULT_1_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(2,4)<=signed(MULT_1_5(2,4)(MULT_SIZE-1) & MULT_1_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(2,4)(MULT_SIZE-1) & MULT_1_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(2,4)<=signed(MULT_2_1(2,4)(MULT_SIZE-1) & MULT_2_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(2,4)(MULT_SIZE-1) & MULT_2_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(2,4)<=signed(MULT_2_3(2,4)(MULT_SIZE-1) & MULT_2_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(2,4)(MULT_SIZE-1) & MULT_2_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(2,4)<=signed(MULT_2_5(2,4)(MULT_SIZE-1) & MULT_2_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(2,4)(MULT_SIZE-1) & MULT_2_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(2,4)<=signed(MULT_3_1(2,4)(MULT_SIZE-1) & MULT_3_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(2,4)(MULT_SIZE-1) & MULT_3_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(2,4)<=signed(MULT_3_3(2,4)(MULT_SIZE-1) & MULT_3_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(2,4)(MULT_SIZE-1) & MULT_3_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(2,4)<=signed(MULT_3_5(2,4)(MULT_SIZE-1) & MULT_3_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(2,4)(MULT_SIZE-1) & MULT_3_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(2,4)<=signed(MULT_4_1(2,4)(MULT_SIZE-1) & MULT_4_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(2,4)(MULT_SIZE-1) & MULT_4_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(2,4)<=signed(MULT_4_3(2,4)(MULT_SIZE-1) & MULT_4_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(2,4)(MULT_SIZE-1) & MULT_4_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(2,4)<=signed(MULT_4_5(2,4)(MULT_SIZE-1) & MULT_4_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(2,4)(MULT_SIZE-1) & MULT_4_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(2,4)<=signed(MULT_5_1(2,4)(MULT_SIZE-1) & MULT_5_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(2,4)(MULT_SIZE-1) & MULT_5_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(2,4)<=signed(MULT_5_3(2,4)(MULT_SIZE-1) & MULT_5_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(2,4)(MULT_SIZE-1) & MULT_5_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(2,4)<=signed(MULT_5_5(2,4)(MULT_SIZE-1) & MULT_5_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(2,4)(MULT_SIZE-1) & MULT_5_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(2,4)<=signed(MULT_6_1(2,4)(MULT_SIZE-1) & MULT_6_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(2,4)(MULT_SIZE-1) & MULT_6_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(2,4)<=signed(MULT_6_3(2,4)(MULT_SIZE-1) & MULT_6_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(2,4)(MULT_SIZE-1) & MULT_6_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(2,4)<=signed(MULT_6_5(2,4)(MULT_SIZE-1) & MULT_6_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(2,4)(MULT_SIZE-1) & MULT_6_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(2,4)<=signed(MULT_7_1(2,4)(MULT_SIZE-1) & MULT_7_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(2,4)(MULT_SIZE-1) & MULT_7_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(2,4)<=signed(MULT_7_3(2,4)(MULT_SIZE-1) & MULT_7_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(2,4)(MULT_SIZE-1) & MULT_7_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(2,4)<=signed(MULT_7_5(2,4)(MULT_SIZE-1) & MULT_7_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(2,4)(MULT_SIZE-1) & MULT_7_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(2,4)<=signed(MULT_8_1(2,4)(MULT_SIZE-1) & MULT_8_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(2,4)(MULT_SIZE-1) & MULT_8_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(2,4)<=signed(MULT_8_3(2,4)(MULT_SIZE-1) & MULT_8_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(2,4)(MULT_SIZE-1) & MULT_8_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(2,4)<=signed(MULT_8_5(2,4)(MULT_SIZE-1) & MULT_8_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(2,4)(MULT_SIZE-1) & MULT_8_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(2,4)<=signed(MULT_9_1(2,4)(MULT_SIZE-1) & MULT_9_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(2,4)(MULT_SIZE-1) & MULT_9_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(2,4)<=signed(MULT_9_3(2,4)(MULT_SIZE-1) & MULT_9_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(2,4)(MULT_SIZE-1) & MULT_9_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(2,4)<=signed(MULT_9_5(2,4)(MULT_SIZE-1) & MULT_9_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(2,4)(MULT_SIZE-1) & MULT_9_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(2,4)<=signed(MULT_10_1(2,4)(MULT_SIZE-1) & MULT_10_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(2,4)(MULT_SIZE-1) & MULT_10_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(2,4)<=signed(MULT_10_3(2,4)(MULT_SIZE-1) & MULT_10_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(2,4)(MULT_SIZE-1) & MULT_10_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(2,4)<=signed(MULT_10_5(2,4)(MULT_SIZE-1) & MULT_10_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(2,4)(MULT_SIZE-1) & MULT_10_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(2,4)<=signed(MULT_11_1(2,4)(MULT_SIZE-1) & MULT_11_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(2,4)(MULT_SIZE-1) & MULT_11_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(2,4)<=signed(MULT_11_3(2,4)(MULT_SIZE-1) & MULT_11_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(2,4)(MULT_SIZE-1) & MULT_11_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(2,4)<=signed(MULT_11_5(2,4)(MULT_SIZE-1) & MULT_11_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(2,4)(MULT_SIZE-1) & MULT_11_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(2,4)<=signed(MULT_12_1(2,4)(MULT_SIZE-1) & MULT_12_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(2,4)(MULT_SIZE-1) & MULT_12_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(2,4)<=signed(MULT_12_3(2,4)(MULT_SIZE-1) & MULT_12_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(2,4)(MULT_SIZE-1) & MULT_12_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(2,4)<=signed(MULT_12_5(2,4)(MULT_SIZE-1) & MULT_12_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(2,4)(MULT_SIZE-1) & MULT_12_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(2,4)<=signed(MULT_13_1(2,4)(MULT_SIZE-1) & MULT_13_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(2,4)(MULT_SIZE-1) & MULT_13_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(2,4)<=signed(MULT_13_3(2,4)(MULT_SIZE-1) & MULT_13_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(2,4)(MULT_SIZE-1) & MULT_13_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(2,4)<=signed(MULT_13_5(2,4)(MULT_SIZE-1) & MULT_13_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(2,4)(MULT_SIZE-1) & MULT_13_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(2,4)<=signed(MULT_14_1(2,4)(MULT_SIZE-1) & MULT_14_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(2,4)(MULT_SIZE-1) & MULT_14_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(2,4)<=signed(MULT_14_3(2,4)(MULT_SIZE-1) & MULT_14_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(2,4)(MULT_SIZE-1) & MULT_14_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(2,4)<=signed(MULT_14_5(2,4)(MULT_SIZE-1) & MULT_14_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(2,4)(MULT_SIZE-1) & MULT_14_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(2,4)<=signed(MULT_15_1(2,4)(MULT_SIZE-1) & MULT_15_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(2,4)(MULT_SIZE-1) & MULT_15_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(2,4)<=signed(MULT_15_3(2,4)(MULT_SIZE-1) & MULT_15_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(2,4)(MULT_SIZE-1) & MULT_15_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(2,4)<=signed(MULT_15_5(2,4)(MULT_SIZE-1) & MULT_15_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(2,4)(MULT_SIZE-1) & MULT_15_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(2,4)<=signed(MULT_16_1(2,4)(MULT_SIZE-1) & MULT_16_1(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(2,4)(MULT_SIZE-1) & MULT_16_2(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(2,4)<=signed(MULT_16_3(2,4)(MULT_SIZE-1) & MULT_16_3(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(2,4)(MULT_SIZE-1) & MULT_16_4(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(2,4)<=signed(MULT_16_5(2,4)(MULT_SIZE-1) & MULT_16_5(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(2,4)(MULT_SIZE-1) & MULT_16_6(2,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(2,4) ------------------

			MULTS_1_1_1(3,0)<=signed(MULT_1_1(3,0)(MULT_SIZE-1) & MULT_1_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(3,0)(MULT_SIZE-1) & MULT_1_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(3,0)<=signed(MULT_1_3(3,0)(MULT_SIZE-1) & MULT_1_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(3,0)(MULT_SIZE-1) & MULT_1_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(3,0)<=signed(MULT_1_5(3,0)(MULT_SIZE-1) & MULT_1_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(3,0)(MULT_SIZE-1) & MULT_1_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(3,0)<=signed(MULT_2_1(3,0)(MULT_SIZE-1) & MULT_2_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(3,0)(MULT_SIZE-1) & MULT_2_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(3,0)<=signed(MULT_2_3(3,0)(MULT_SIZE-1) & MULT_2_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(3,0)(MULT_SIZE-1) & MULT_2_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(3,0)<=signed(MULT_2_5(3,0)(MULT_SIZE-1) & MULT_2_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(3,0)(MULT_SIZE-1) & MULT_2_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(3,0)<=signed(MULT_3_1(3,0)(MULT_SIZE-1) & MULT_3_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(3,0)(MULT_SIZE-1) & MULT_3_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(3,0)<=signed(MULT_3_3(3,0)(MULT_SIZE-1) & MULT_3_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(3,0)(MULT_SIZE-1) & MULT_3_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(3,0)<=signed(MULT_3_5(3,0)(MULT_SIZE-1) & MULT_3_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(3,0)(MULT_SIZE-1) & MULT_3_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(3,0)<=signed(MULT_4_1(3,0)(MULT_SIZE-1) & MULT_4_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(3,0)(MULT_SIZE-1) & MULT_4_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(3,0)<=signed(MULT_4_3(3,0)(MULT_SIZE-1) & MULT_4_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(3,0)(MULT_SIZE-1) & MULT_4_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(3,0)<=signed(MULT_4_5(3,0)(MULT_SIZE-1) & MULT_4_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(3,0)(MULT_SIZE-1) & MULT_4_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(3,0)<=signed(MULT_5_1(3,0)(MULT_SIZE-1) & MULT_5_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(3,0)(MULT_SIZE-1) & MULT_5_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(3,0)<=signed(MULT_5_3(3,0)(MULT_SIZE-1) & MULT_5_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(3,0)(MULT_SIZE-1) & MULT_5_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(3,0)<=signed(MULT_5_5(3,0)(MULT_SIZE-1) & MULT_5_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(3,0)(MULT_SIZE-1) & MULT_5_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(3,0)<=signed(MULT_6_1(3,0)(MULT_SIZE-1) & MULT_6_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(3,0)(MULT_SIZE-1) & MULT_6_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(3,0)<=signed(MULT_6_3(3,0)(MULT_SIZE-1) & MULT_6_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(3,0)(MULT_SIZE-1) & MULT_6_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(3,0)<=signed(MULT_6_5(3,0)(MULT_SIZE-1) & MULT_6_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(3,0)(MULT_SIZE-1) & MULT_6_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(3,0)<=signed(MULT_7_1(3,0)(MULT_SIZE-1) & MULT_7_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(3,0)(MULT_SIZE-1) & MULT_7_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(3,0)<=signed(MULT_7_3(3,0)(MULT_SIZE-1) & MULT_7_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(3,0)(MULT_SIZE-1) & MULT_7_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(3,0)<=signed(MULT_7_5(3,0)(MULT_SIZE-1) & MULT_7_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(3,0)(MULT_SIZE-1) & MULT_7_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(3,0)<=signed(MULT_8_1(3,0)(MULT_SIZE-1) & MULT_8_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(3,0)(MULT_SIZE-1) & MULT_8_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(3,0)<=signed(MULT_8_3(3,0)(MULT_SIZE-1) & MULT_8_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(3,0)(MULT_SIZE-1) & MULT_8_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(3,0)<=signed(MULT_8_5(3,0)(MULT_SIZE-1) & MULT_8_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(3,0)(MULT_SIZE-1) & MULT_8_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(3,0)<=signed(MULT_9_1(3,0)(MULT_SIZE-1) & MULT_9_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(3,0)(MULT_SIZE-1) & MULT_9_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(3,0)<=signed(MULT_9_3(3,0)(MULT_SIZE-1) & MULT_9_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(3,0)(MULT_SIZE-1) & MULT_9_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(3,0)<=signed(MULT_9_5(3,0)(MULT_SIZE-1) & MULT_9_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(3,0)(MULT_SIZE-1) & MULT_9_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(3,0)<=signed(MULT_10_1(3,0)(MULT_SIZE-1) & MULT_10_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(3,0)(MULT_SIZE-1) & MULT_10_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(3,0)<=signed(MULT_10_3(3,0)(MULT_SIZE-1) & MULT_10_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(3,0)(MULT_SIZE-1) & MULT_10_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(3,0)<=signed(MULT_10_5(3,0)(MULT_SIZE-1) & MULT_10_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(3,0)(MULT_SIZE-1) & MULT_10_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(3,0)<=signed(MULT_11_1(3,0)(MULT_SIZE-1) & MULT_11_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(3,0)(MULT_SIZE-1) & MULT_11_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(3,0)<=signed(MULT_11_3(3,0)(MULT_SIZE-1) & MULT_11_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(3,0)(MULT_SIZE-1) & MULT_11_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(3,0)<=signed(MULT_11_5(3,0)(MULT_SIZE-1) & MULT_11_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(3,0)(MULT_SIZE-1) & MULT_11_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(3,0)<=signed(MULT_12_1(3,0)(MULT_SIZE-1) & MULT_12_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(3,0)(MULT_SIZE-1) & MULT_12_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(3,0)<=signed(MULT_12_3(3,0)(MULT_SIZE-1) & MULT_12_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(3,0)(MULT_SIZE-1) & MULT_12_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(3,0)<=signed(MULT_12_5(3,0)(MULT_SIZE-1) & MULT_12_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(3,0)(MULT_SIZE-1) & MULT_12_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(3,0)<=signed(MULT_13_1(3,0)(MULT_SIZE-1) & MULT_13_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(3,0)(MULT_SIZE-1) & MULT_13_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(3,0)<=signed(MULT_13_3(3,0)(MULT_SIZE-1) & MULT_13_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(3,0)(MULT_SIZE-1) & MULT_13_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(3,0)<=signed(MULT_13_5(3,0)(MULT_SIZE-1) & MULT_13_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(3,0)(MULT_SIZE-1) & MULT_13_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(3,0)<=signed(MULT_14_1(3,0)(MULT_SIZE-1) & MULT_14_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(3,0)(MULT_SIZE-1) & MULT_14_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(3,0)<=signed(MULT_14_3(3,0)(MULT_SIZE-1) & MULT_14_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(3,0)(MULT_SIZE-1) & MULT_14_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(3,0)<=signed(MULT_14_5(3,0)(MULT_SIZE-1) & MULT_14_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(3,0)(MULT_SIZE-1) & MULT_14_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(3,0)<=signed(MULT_15_1(3,0)(MULT_SIZE-1) & MULT_15_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(3,0)(MULT_SIZE-1) & MULT_15_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(3,0)<=signed(MULT_15_3(3,0)(MULT_SIZE-1) & MULT_15_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(3,0)(MULT_SIZE-1) & MULT_15_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(3,0)<=signed(MULT_15_5(3,0)(MULT_SIZE-1) & MULT_15_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(3,0)(MULT_SIZE-1) & MULT_15_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(3,0)<=signed(MULT_16_1(3,0)(MULT_SIZE-1) & MULT_16_1(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(3,0)(MULT_SIZE-1) & MULT_16_2(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(3,0)<=signed(MULT_16_3(3,0)(MULT_SIZE-1) & MULT_16_3(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(3,0)(MULT_SIZE-1) & MULT_16_4(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(3,0)<=signed(MULT_16_5(3,0)(MULT_SIZE-1) & MULT_16_5(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(3,0)(MULT_SIZE-1) & MULT_16_6(3,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(3,0) ------------------

			MULTS_1_1_1(3,1)<=signed(MULT_1_1(3,1)(MULT_SIZE-1) & MULT_1_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(3,1)(MULT_SIZE-1) & MULT_1_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(3,1)<=signed(MULT_1_3(3,1)(MULT_SIZE-1) & MULT_1_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(3,1)(MULT_SIZE-1) & MULT_1_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(3,1)<=signed(MULT_1_5(3,1)(MULT_SIZE-1) & MULT_1_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(3,1)(MULT_SIZE-1) & MULT_1_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(3,1)<=signed(MULT_2_1(3,1)(MULT_SIZE-1) & MULT_2_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(3,1)(MULT_SIZE-1) & MULT_2_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(3,1)<=signed(MULT_2_3(3,1)(MULT_SIZE-1) & MULT_2_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(3,1)(MULT_SIZE-1) & MULT_2_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(3,1)<=signed(MULT_2_5(3,1)(MULT_SIZE-1) & MULT_2_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(3,1)(MULT_SIZE-1) & MULT_2_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(3,1)<=signed(MULT_3_1(3,1)(MULT_SIZE-1) & MULT_3_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(3,1)(MULT_SIZE-1) & MULT_3_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(3,1)<=signed(MULT_3_3(3,1)(MULT_SIZE-1) & MULT_3_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(3,1)(MULT_SIZE-1) & MULT_3_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(3,1)<=signed(MULT_3_5(3,1)(MULT_SIZE-1) & MULT_3_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(3,1)(MULT_SIZE-1) & MULT_3_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(3,1)<=signed(MULT_4_1(3,1)(MULT_SIZE-1) & MULT_4_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(3,1)(MULT_SIZE-1) & MULT_4_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(3,1)<=signed(MULT_4_3(3,1)(MULT_SIZE-1) & MULT_4_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(3,1)(MULT_SIZE-1) & MULT_4_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(3,1)<=signed(MULT_4_5(3,1)(MULT_SIZE-1) & MULT_4_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(3,1)(MULT_SIZE-1) & MULT_4_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(3,1)<=signed(MULT_5_1(3,1)(MULT_SIZE-1) & MULT_5_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(3,1)(MULT_SIZE-1) & MULT_5_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(3,1)<=signed(MULT_5_3(3,1)(MULT_SIZE-1) & MULT_5_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(3,1)(MULT_SIZE-1) & MULT_5_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(3,1)<=signed(MULT_5_5(3,1)(MULT_SIZE-1) & MULT_5_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(3,1)(MULT_SIZE-1) & MULT_5_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(3,1)<=signed(MULT_6_1(3,1)(MULT_SIZE-1) & MULT_6_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(3,1)(MULT_SIZE-1) & MULT_6_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(3,1)<=signed(MULT_6_3(3,1)(MULT_SIZE-1) & MULT_6_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(3,1)(MULT_SIZE-1) & MULT_6_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(3,1)<=signed(MULT_6_5(3,1)(MULT_SIZE-1) & MULT_6_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(3,1)(MULT_SIZE-1) & MULT_6_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(3,1)<=signed(MULT_7_1(3,1)(MULT_SIZE-1) & MULT_7_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(3,1)(MULT_SIZE-1) & MULT_7_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(3,1)<=signed(MULT_7_3(3,1)(MULT_SIZE-1) & MULT_7_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(3,1)(MULT_SIZE-1) & MULT_7_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(3,1)<=signed(MULT_7_5(3,1)(MULT_SIZE-1) & MULT_7_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(3,1)(MULT_SIZE-1) & MULT_7_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(3,1)<=signed(MULT_8_1(3,1)(MULT_SIZE-1) & MULT_8_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(3,1)(MULT_SIZE-1) & MULT_8_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(3,1)<=signed(MULT_8_3(3,1)(MULT_SIZE-1) & MULT_8_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(3,1)(MULT_SIZE-1) & MULT_8_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(3,1)<=signed(MULT_8_5(3,1)(MULT_SIZE-1) & MULT_8_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(3,1)(MULT_SIZE-1) & MULT_8_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(3,1)<=signed(MULT_9_1(3,1)(MULT_SIZE-1) & MULT_9_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(3,1)(MULT_SIZE-1) & MULT_9_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(3,1)<=signed(MULT_9_3(3,1)(MULT_SIZE-1) & MULT_9_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(3,1)(MULT_SIZE-1) & MULT_9_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(3,1)<=signed(MULT_9_5(3,1)(MULT_SIZE-1) & MULT_9_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(3,1)(MULT_SIZE-1) & MULT_9_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(3,1)<=signed(MULT_10_1(3,1)(MULT_SIZE-1) & MULT_10_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(3,1)(MULT_SIZE-1) & MULT_10_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(3,1)<=signed(MULT_10_3(3,1)(MULT_SIZE-1) & MULT_10_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(3,1)(MULT_SIZE-1) & MULT_10_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(3,1)<=signed(MULT_10_5(3,1)(MULT_SIZE-1) & MULT_10_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(3,1)(MULT_SIZE-1) & MULT_10_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(3,1)<=signed(MULT_11_1(3,1)(MULT_SIZE-1) & MULT_11_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(3,1)(MULT_SIZE-1) & MULT_11_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(3,1)<=signed(MULT_11_3(3,1)(MULT_SIZE-1) & MULT_11_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(3,1)(MULT_SIZE-1) & MULT_11_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(3,1)<=signed(MULT_11_5(3,1)(MULT_SIZE-1) & MULT_11_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(3,1)(MULT_SIZE-1) & MULT_11_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(3,1)<=signed(MULT_12_1(3,1)(MULT_SIZE-1) & MULT_12_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(3,1)(MULT_SIZE-1) & MULT_12_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(3,1)<=signed(MULT_12_3(3,1)(MULT_SIZE-1) & MULT_12_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(3,1)(MULT_SIZE-1) & MULT_12_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(3,1)<=signed(MULT_12_5(3,1)(MULT_SIZE-1) & MULT_12_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(3,1)(MULT_SIZE-1) & MULT_12_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(3,1)<=signed(MULT_13_1(3,1)(MULT_SIZE-1) & MULT_13_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(3,1)(MULT_SIZE-1) & MULT_13_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(3,1)<=signed(MULT_13_3(3,1)(MULT_SIZE-1) & MULT_13_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(3,1)(MULT_SIZE-1) & MULT_13_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(3,1)<=signed(MULT_13_5(3,1)(MULT_SIZE-1) & MULT_13_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(3,1)(MULT_SIZE-1) & MULT_13_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(3,1)<=signed(MULT_14_1(3,1)(MULT_SIZE-1) & MULT_14_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(3,1)(MULT_SIZE-1) & MULT_14_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(3,1)<=signed(MULT_14_3(3,1)(MULT_SIZE-1) & MULT_14_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(3,1)(MULT_SIZE-1) & MULT_14_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(3,1)<=signed(MULT_14_5(3,1)(MULT_SIZE-1) & MULT_14_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(3,1)(MULT_SIZE-1) & MULT_14_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(3,1)<=signed(MULT_15_1(3,1)(MULT_SIZE-1) & MULT_15_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(3,1)(MULT_SIZE-1) & MULT_15_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(3,1)<=signed(MULT_15_3(3,1)(MULT_SIZE-1) & MULT_15_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(3,1)(MULT_SIZE-1) & MULT_15_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(3,1)<=signed(MULT_15_5(3,1)(MULT_SIZE-1) & MULT_15_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(3,1)(MULT_SIZE-1) & MULT_15_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(3,1)<=signed(MULT_16_1(3,1)(MULT_SIZE-1) & MULT_16_1(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(3,1)(MULT_SIZE-1) & MULT_16_2(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(3,1)<=signed(MULT_16_3(3,1)(MULT_SIZE-1) & MULT_16_3(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(3,1)(MULT_SIZE-1) & MULT_16_4(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(3,1)<=signed(MULT_16_5(3,1)(MULT_SIZE-1) & MULT_16_5(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(3,1)(MULT_SIZE-1) & MULT_16_6(3,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(3,1) ------------------

			MULTS_1_1_1(3,2)<=signed(MULT_1_1(3,2)(MULT_SIZE-1) & MULT_1_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(3,2)(MULT_SIZE-1) & MULT_1_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(3,2)<=signed(MULT_1_3(3,2)(MULT_SIZE-1) & MULT_1_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(3,2)(MULT_SIZE-1) & MULT_1_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(3,2)<=signed(MULT_1_5(3,2)(MULT_SIZE-1) & MULT_1_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(3,2)(MULT_SIZE-1) & MULT_1_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(3,2)<=signed(MULT_2_1(3,2)(MULT_SIZE-1) & MULT_2_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(3,2)(MULT_SIZE-1) & MULT_2_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(3,2)<=signed(MULT_2_3(3,2)(MULT_SIZE-1) & MULT_2_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(3,2)(MULT_SIZE-1) & MULT_2_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(3,2)<=signed(MULT_2_5(3,2)(MULT_SIZE-1) & MULT_2_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(3,2)(MULT_SIZE-1) & MULT_2_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(3,2)<=signed(MULT_3_1(3,2)(MULT_SIZE-1) & MULT_3_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(3,2)(MULT_SIZE-1) & MULT_3_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(3,2)<=signed(MULT_3_3(3,2)(MULT_SIZE-1) & MULT_3_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(3,2)(MULT_SIZE-1) & MULT_3_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(3,2)<=signed(MULT_3_5(3,2)(MULT_SIZE-1) & MULT_3_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(3,2)(MULT_SIZE-1) & MULT_3_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(3,2)<=signed(MULT_4_1(3,2)(MULT_SIZE-1) & MULT_4_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(3,2)(MULT_SIZE-1) & MULT_4_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(3,2)<=signed(MULT_4_3(3,2)(MULT_SIZE-1) & MULT_4_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(3,2)(MULT_SIZE-1) & MULT_4_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(3,2)<=signed(MULT_4_5(3,2)(MULT_SIZE-1) & MULT_4_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(3,2)(MULT_SIZE-1) & MULT_4_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(3,2)<=signed(MULT_5_1(3,2)(MULT_SIZE-1) & MULT_5_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(3,2)(MULT_SIZE-1) & MULT_5_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(3,2)<=signed(MULT_5_3(3,2)(MULT_SIZE-1) & MULT_5_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(3,2)(MULT_SIZE-1) & MULT_5_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(3,2)<=signed(MULT_5_5(3,2)(MULT_SIZE-1) & MULT_5_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(3,2)(MULT_SIZE-1) & MULT_5_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(3,2)<=signed(MULT_6_1(3,2)(MULT_SIZE-1) & MULT_6_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(3,2)(MULT_SIZE-1) & MULT_6_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(3,2)<=signed(MULT_6_3(3,2)(MULT_SIZE-1) & MULT_6_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(3,2)(MULT_SIZE-1) & MULT_6_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(3,2)<=signed(MULT_6_5(3,2)(MULT_SIZE-1) & MULT_6_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(3,2)(MULT_SIZE-1) & MULT_6_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(3,2)<=signed(MULT_7_1(3,2)(MULT_SIZE-1) & MULT_7_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(3,2)(MULT_SIZE-1) & MULT_7_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(3,2)<=signed(MULT_7_3(3,2)(MULT_SIZE-1) & MULT_7_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(3,2)(MULT_SIZE-1) & MULT_7_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(3,2)<=signed(MULT_7_5(3,2)(MULT_SIZE-1) & MULT_7_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(3,2)(MULT_SIZE-1) & MULT_7_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(3,2)<=signed(MULT_8_1(3,2)(MULT_SIZE-1) & MULT_8_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(3,2)(MULT_SIZE-1) & MULT_8_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(3,2)<=signed(MULT_8_3(3,2)(MULT_SIZE-1) & MULT_8_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(3,2)(MULT_SIZE-1) & MULT_8_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(3,2)<=signed(MULT_8_5(3,2)(MULT_SIZE-1) & MULT_8_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(3,2)(MULT_SIZE-1) & MULT_8_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(3,2)<=signed(MULT_9_1(3,2)(MULT_SIZE-1) & MULT_9_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(3,2)(MULT_SIZE-1) & MULT_9_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(3,2)<=signed(MULT_9_3(3,2)(MULT_SIZE-1) & MULT_9_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(3,2)(MULT_SIZE-1) & MULT_9_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(3,2)<=signed(MULT_9_5(3,2)(MULT_SIZE-1) & MULT_9_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(3,2)(MULT_SIZE-1) & MULT_9_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(3,2)<=signed(MULT_10_1(3,2)(MULT_SIZE-1) & MULT_10_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(3,2)(MULT_SIZE-1) & MULT_10_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(3,2)<=signed(MULT_10_3(3,2)(MULT_SIZE-1) & MULT_10_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(3,2)(MULT_SIZE-1) & MULT_10_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(3,2)<=signed(MULT_10_5(3,2)(MULT_SIZE-1) & MULT_10_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(3,2)(MULT_SIZE-1) & MULT_10_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(3,2)<=signed(MULT_11_1(3,2)(MULT_SIZE-1) & MULT_11_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(3,2)(MULT_SIZE-1) & MULT_11_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(3,2)<=signed(MULT_11_3(3,2)(MULT_SIZE-1) & MULT_11_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(3,2)(MULT_SIZE-1) & MULT_11_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(3,2)<=signed(MULT_11_5(3,2)(MULT_SIZE-1) & MULT_11_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(3,2)(MULT_SIZE-1) & MULT_11_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(3,2)<=signed(MULT_12_1(3,2)(MULT_SIZE-1) & MULT_12_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(3,2)(MULT_SIZE-1) & MULT_12_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(3,2)<=signed(MULT_12_3(3,2)(MULT_SIZE-1) & MULT_12_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(3,2)(MULT_SIZE-1) & MULT_12_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(3,2)<=signed(MULT_12_5(3,2)(MULT_SIZE-1) & MULT_12_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(3,2)(MULT_SIZE-1) & MULT_12_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(3,2)<=signed(MULT_13_1(3,2)(MULT_SIZE-1) & MULT_13_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(3,2)(MULT_SIZE-1) & MULT_13_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(3,2)<=signed(MULT_13_3(3,2)(MULT_SIZE-1) & MULT_13_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(3,2)(MULT_SIZE-1) & MULT_13_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(3,2)<=signed(MULT_13_5(3,2)(MULT_SIZE-1) & MULT_13_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(3,2)(MULT_SIZE-1) & MULT_13_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(3,2)<=signed(MULT_14_1(3,2)(MULT_SIZE-1) & MULT_14_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(3,2)(MULT_SIZE-1) & MULT_14_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(3,2)<=signed(MULT_14_3(3,2)(MULT_SIZE-1) & MULT_14_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(3,2)(MULT_SIZE-1) & MULT_14_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(3,2)<=signed(MULT_14_5(3,2)(MULT_SIZE-1) & MULT_14_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(3,2)(MULT_SIZE-1) & MULT_14_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(3,2)<=signed(MULT_15_1(3,2)(MULT_SIZE-1) & MULT_15_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(3,2)(MULT_SIZE-1) & MULT_15_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(3,2)<=signed(MULT_15_3(3,2)(MULT_SIZE-1) & MULT_15_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(3,2)(MULT_SIZE-1) & MULT_15_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(3,2)<=signed(MULT_15_5(3,2)(MULT_SIZE-1) & MULT_15_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(3,2)(MULT_SIZE-1) & MULT_15_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(3,2)<=signed(MULT_16_1(3,2)(MULT_SIZE-1) & MULT_16_1(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(3,2)(MULT_SIZE-1) & MULT_16_2(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(3,2)<=signed(MULT_16_3(3,2)(MULT_SIZE-1) & MULT_16_3(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(3,2)(MULT_SIZE-1) & MULT_16_4(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(3,2)<=signed(MULT_16_5(3,2)(MULT_SIZE-1) & MULT_16_5(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(3,2)(MULT_SIZE-1) & MULT_16_6(3,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(3,2) ------------------

			MULTS_1_1_1(3,3)<=signed(MULT_1_1(3,3)(MULT_SIZE-1) & MULT_1_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(3,3)(MULT_SIZE-1) & MULT_1_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(3,3)<=signed(MULT_1_3(3,3)(MULT_SIZE-1) & MULT_1_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(3,3)(MULT_SIZE-1) & MULT_1_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(3,3)<=signed(MULT_1_5(3,3)(MULT_SIZE-1) & MULT_1_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(3,3)(MULT_SIZE-1) & MULT_1_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(3,3)<=signed(MULT_2_1(3,3)(MULT_SIZE-1) & MULT_2_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(3,3)(MULT_SIZE-1) & MULT_2_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(3,3)<=signed(MULT_2_3(3,3)(MULT_SIZE-1) & MULT_2_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(3,3)(MULT_SIZE-1) & MULT_2_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(3,3)<=signed(MULT_2_5(3,3)(MULT_SIZE-1) & MULT_2_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(3,3)(MULT_SIZE-1) & MULT_2_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(3,3)<=signed(MULT_3_1(3,3)(MULT_SIZE-1) & MULT_3_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(3,3)(MULT_SIZE-1) & MULT_3_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(3,3)<=signed(MULT_3_3(3,3)(MULT_SIZE-1) & MULT_3_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(3,3)(MULT_SIZE-1) & MULT_3_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(3,3)<=signed(MULT_3_5(3,3)(MULT_SIZE-1) & MULT_3_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(3,3)(MULT_SIZE-1) & MULT_3_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(3,3)<=signed(MULT_4_1(3,3)(MULT_SIZE-1) & MULT_4_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(3,3)(MULT_SIZE-1) & MULT_4_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(3,3)<=signed(MULT_4_3(3,3)(MULT_SIZE-1) & MULT_4_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(3,3)(MULT_SIZE-1) & MULT_4_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(3,3)<=signed(MULT_4_5(3,3)(MULT_SIZE-1) & MULT_4_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(3,3)(MULT_SIZE-1) & MULT_4_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(3,3)<=signed(MULT_5_1(3,3)(MULT_SIZE-1) & MULT_5_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(3,3)(MULT_SIZE-1) & MULT_5_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(3,3)<=signed(MULT_5_3(3,3)(MULT_SIZE-1) & MULT_5_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(3,3)(MULT_SIZE-1) & MULT_5_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(3,3)<=signed(MULT_5_5(3,3)(MULT_SIZE-1) & MULT_5_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(3,3)(MULT_SIZE-1) & MULT_5_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(3,3)<=signed(MULT_6_1(3,3)(MULT_SIZE-1) & MULT_6_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(3,3)(MULT_SIZE-1) & MULT_6_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(3,3)<=signed(MULT_6_3(3,3)(MULT_SIZE-1) & MULT_6_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(3,3)(MULT_SIZE-1) & MULT_6_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(3,3)<=signed(MULT_6_5(3,3)(MULT_SIZE-1) & MULT_6_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(3,3)(MULT_SIZE-1) & MULT_6_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(3,3)<=signed(MULT_7_1(3,3)(MULT_SIZE-1) & MULT_7_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(3,3)(MULT_SIZE-1) & MULT_7_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(3,3)<=signed(MULT_7_3(3,3)(MULT_SIZE-1) & MULT_7_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(3,3)(MULT_SIZE-1) & MULT_7_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(3,3)<=signed(MULT_7_5(3,3)(MULT_SIZE-1) & MULT_7_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(3,3)(MULT_SIZE-1) & MULT_7_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(3,3)<=signed(MULT_8_1(3,3)(MULT_SIZE-1) & MULT_8_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(3,3)(MULT_SIZE-1) & MULT_8_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(3,3)<=signed(MULT_8_3(3,3)(MULT_SIZE-1) & MULT_8_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(3,3)(MULT_SIZE-1) & MULT_8_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(3,3)<=signed(MULT_8_5(3,3)(MULT_SIZE-1) & MULT_8_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(3,3)(MULT_SIZE-1) & MULT_8_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(3,3)<=signed(MULT_9_1(3,3)(MULT_SIZE-1) & MULT_9_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(3,3)(MULT_SIZE-1) & MULT_9_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(3,3)<=signed(MULT_9_3(3,3)(MULT_SIZE-1) & MULT_9_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(3,3)(MULT_SIZE-1) & MULT_9_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(3,3)<=signed(MULT_9_5(3,3)(MULT_SIZE-1) & MULT_9_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(3,3)(MULT_SIZE-1) & MULT_9_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(3,3)<=signed(MULT_10_1(3,3)(MULT_SIZE-1) & MULT_10_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(3,3)(MULT_SIZE-1) & MULT_10_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(3,3)<=signed(MULT_10_3(3,3)(MULT_SIZE-1) & MULT_10_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(3,3)(MULT_SIZE-1) & MULT_10_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(3,3)<=signed(MULT_10_5(3,3)(MULT_SIZE-1) & MULT_10_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(3,3)(MULT_SIZE-1) & MULT_10_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(3,3)<=signed(MULT_11_1(3,3)(MULT_SIZE-1) & MULT_11_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(3,3)(MULT_SIZE-1) & MULT_11_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(3,3)<=signed(MULT_11_3(3,3)(MULT_SIZE-1) & MULT_11_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(3,3)(MULT_SIZE-1) & MULT_11_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(3,3)<=signed(MULT_11_5(3,3)(MULT_SIZE-1) & MULT_11_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(3,3)(MULT_SIZE-1) & MULT_11_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(3,3)<=signed(MULT_12_1(3,3)(MULT_SIZE-1) & MULT_12_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(3,3)(MULT_SIZE-1) & MULT_12_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(3,3)<=signed(MULT_12_3(3,3)(MULT_SIZE-1) & MULT_12_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(3,3)(MULT_SIZE-1) & MULT_12_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(3,3)<=signed(MULT_12_5(3,3)(MULT_SIZE-1) & MULT_12_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(3,3)(MULT_SIZE-1) & MULT_12_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(3,3)<=signed(MULT_13_1(3,3)(MULT_SIZE-1) & MULT_13_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(3,3)(MULT_SIZE-1) & MULT_13_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(3,3)<=signed(MULT_13_3(3,3)(MULT_SIZE-1) & MULT_13_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(3,3)(MULT_SIZE-1) & MULT_13_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(3,3)<=signed(MULT_13_5(3,3)(MULT_SIZE-1) & MULT_13_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(3,3)(MULT_SIZE-1) & MULT_13_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(3,3)<=signed(MULT_14_1(3,3)(MULT_SIZE-1) & MULT_14_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(3,3)(MULT_SIZE-1) & MULT_14_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(3,3)<=signed(MULT_14_3(3,3)(MULT_SIZE-1) & MULT_14_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(3,3)(MULT_SIZE-1) & MULT_14_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(3,3)<=signed(MULT_14_5(3,3)(MULT_SIZE-1) & MULT_14_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(3,3)(MULT_SIZE-1) & MULT_14_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(3,3)<=signed(MULT_15_1(3,3)(MULT_SIZE-1) & MULT_15_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(3,3)(MULT_SIZE-1) & MULT_15_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(3,3)<=signed(MULT_15_3(3,3)(MULT_SIZE-1) & MULT_15_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(3,3)(MULT_SIZE-1) & MULT_15_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(3,3)<=signed(MULT_15_5(3,3)(MULT_SIZE-1) & MULT_15_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(3,3)(MULT_SIZE-1) & MULT_15_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(3,3)<=signed(MULT_16_1(3,3)(MULT_SIZE-1) & MULT_16_1(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(3,3)(MULT_SIZE-1) & MULT_16_2(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(3,3)<=signed(MULT_16_3(3,3)(MULT_SIZE-1) & MULT_16_3(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(3,3)(MULT_SIZE-1) & MULT_16_4(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(3,3)<=signed(MULT_16_5(3,3)(MULT_SIZE-1) & MULT_16_5(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(3,3)(MULT_SIZE-1) & MULT_16_6(3,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(3,3) ------------------

			MULTS_1_1_1(3,4)<=signed(MULT_1_1(3,4)(MULT_SIZE-1) & MULT_1_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(3,4)(MULT_SIZE-1) & MULT_1_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(3,4)<=signed(MULT_1_3(3,4)(MULT_SIZE-1) & MULT_1_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(3,4)(MULT_SIZE-1) & MULT_1_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(3,4)<=signed(MULT_1_5(3,4)(MULT_SIZE-1) & MULT_1_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(3,4)(MULT_SIZE-1) & MULT_1_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(3,4)<=signed(MULT_2_1(3,4)(MULT_SIZE-1) & MULT_2_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(3,4)(MULT_SIZE-1) & MULT_2_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(3,4)<=signed(MULT_2_3(3,4)(MULT_SIZE-1) & MULT_2_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(3,4)(MULT_SIZE-1) & MULT_2_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(3,4)<=signed(MULT_2_5(3,4)(MULT_SIZE-1) & MULT_2_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(3,4)(MULT_SIZE-1) & MULT_2_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(3,4)<=signed(MULT_3_1(3,4)(MULT_SIZE-1) & MULT_3_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(3,4)(MULT_SIZE-1) & MULT_3_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(3,4)<=signed(MULT_3_3(3,4)(MULT_SIZE-1) & MULT_3_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(3,4)(MULT_SIZE-1) & MULT_3_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(3,4)<=signed(MULT_3_5(3,4)(MULT_SIZE-1) & MULT_3_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(3,4)(MULT_SIZE-1) & MULT_3_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(3,4)<=signed(MULT_4_1(3,4)(MULT_SIZE-1) & MULT_4_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(3,4)(MULT_SIZE-1) & MULT_4_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(3,4)<=signed(MULT_4_3(3,4)(MULT_SIZE-1) & MULT_4_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(3,4)(MULT_SIZE-1) & MULT_4_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(3,4)<=signed(MULT_4_5(3,4)(MULT_SIZE-1) & MULT_4_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(3,4)(MULT_SIZE-1) & MULT_4_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(3,4)<=signed(MULT_5_1(3,4)(MULT_SIZE-1) & MULT_5_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(3,4)(MULT_SIZE-1) & MULT_5_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(3,4)<=signed(MULT_5_3(3,4)(MULT_SIZE-1) & MULT_5_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(3,4)(MULT_SIZE-1) & MULT_5_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(3,4)<=signed(MULT_5_5(3,4)(MULT_SIZE-1) & MULT_5_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(3,4)(MULT_SIZE-1) & MULT_5_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(3,4)<=signed(MULT_6_1(3,4)(MULT_SIZE-1) & MULT_6_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(3,4)(MULT_SIZE-1) & MULT_6_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(3,4)<=signed(MULT_6_3(3,4)(MULT_SIZE-1) & MULT_6_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(3,4)(MULT_SIZE-1) & MULT_6_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(3,4)<=signed(MULT_6_5(3,4)(MULT_SIZE-1) & MULT_6_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(3,4)(MULT_SIZE-1) & MULT_6_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(3,4)<=signed(MULT_7_1(3,4)(MULT_SIZE-1) & MULT_7_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(3,4)(MULT_SIZE-1) & MULT_7_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(3,4)<=signed(MULT_7_3(3,4)(MULT_SIZE-1) & MULT_7_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(3,4)(MULT_SIZE-1) & MULT_7_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(3,4)<=signed(MULT_7_5(3,4)(MULT_SIZE-1) & MULT_7_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(3,4)(MULT_SIZE-1) & MULT_7_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(3,4)<=signed(MULT_8_1(3,4)(MULT_SIZE-1) & MULT_8_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(3,4)(MULT_SIZE-1) & MULT_8_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(3,4)<=signed(MULT_8_3(3,4)(MULT_SIZE-1) & MULT_8_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(3,4)(MULT_SIZE-1) & MULT_8_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(3,4)<=signed(MULT_8_5(3,4)(MULT_SIZE-1) & MULT_8_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(3,4)(MULT_SIZE-1) & MULT_8_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(3,4)<=signed(MULT_9_1(3,4)(MULT_SIZE-1) & MULT_9_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(3,4)(MULT_SIZE-1) & MULT_9_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(3,4)<=signed(MULT_9_3(3,4)(MULT_SIZE-1) & MULT_9_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(3,4)(MULT_SIZE-1) & MULT_9_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(3,4)<=signed(MULT_9_5(3,4)(MULT_SIZE-1) & MULT_9_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(3,4)(MULT_SIZE-1) & MULT_9_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(3,4)<=signed(MULT_10_1(3,4)(MULT_SIZE-1) & MULT_10_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(3,4)(MULT_SIZE-1) & MULT_10_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(3,4)<=signed(MULT_10_3(3,4)(MULT_SIZE-1) & MULT_10_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(3,4)(MULT_SIZE-1) & MULT_10_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(3,4)<=signed(MULT_10_5(3,4)(MULT_SIZE-1) & MULT_10_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(3,4)(MULT_SIZE-1) & MULT_10_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(3,4)<=signed(MULT_11_1(3,4)(MULT_SIZE-1) & MULT_11_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(3,4)(MULT_SIZE-1) & MULT_11_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(3,4)<=signed(MULT_11_3(3,4)(MULT_SIZE-1) & MULT_11_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(3,4)(MULT_SIZE-1) & MULT_11_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(3,4)<=signed(MULT_11_5(3,4)(MULT_SIZE-1) & MULT_11_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(3,4)(MULT_SIZE-1) & MULT_11_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(3,4)<=signed(MULT_12_1(3,4)(MULT_SIZE-1) & MULT_12_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(3,4)(MULT_SIZE-1) & MULT_12_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(3,4)<=signed(MULT_12_3(3,4)(MULT_SIZE-1) & MULT_12_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(3,4)(MULT_SIZE-1) & MULT_12_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(3,4)<=signed(MULT_12_5(3,4)(MULT_SIZE-1) & MULT_12_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(3,4)(MULT_SIZE-1) & MULT_12_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(3,4)<=signed(MULT_13_1(3,4)(MULT_SIZE-1) & MULT_13_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(3,4)(MULT_SIZE-1) & MULT_13_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(3,4)<=signed(MULT_13_3(3,4)(MULT_SIZE-1) & MULT_13_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(3,4)(MULT_SIZE-1) & MULT_13_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(3,4)<=signed(MULT_13_5(3,4)(MULT_SIZE-1) & MULT_13_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(3,4)(MULT_SIZE-1) & MULT_13_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(3,4)<=signed(MULT_14_1(3,4)(MULT_SIZE-1) & MULT_14_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(3,4)(MULT_SIZE-1) & MULT_14_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(3,4)<=signed(MULT_14_3(3,4)(MULT_SIZE-1) & MULT_14_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(3,4)(MULT_SIZE-1) & MULT_14_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(3,4)<=signed(MULT_14_5(3,4)(MULT_SIZE-1) & MULT_14_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(3,4)(MULT_SIZE-1) & MULT_14_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(3,4)<=signed(MULT_15_1(3,4)(MULT_SIZE-1) & MULT_15_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(3,4)(MULT_SIZE-1) & MULT_15_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(3,4)<=signed(MULT_15_3(3,4)(MULT_SIZE-1) & MULT_15_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(3,4)(MULT_SIZE-1) & MULT_15_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(3,4)<=signed(MULT_15_5(3,4)(MULT_SIZE-1) & MULT_15_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(3,4)(MULT_SIZE-1) & MULT_15_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(3,4)<=signed(MULT_16_1(3,4)(MULT_SIZE-1) & MULT_16_1(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(3,4)(MULT_SIZE-1) & MULT_16_2(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(3,4)<=signed(MULT_16_3(3,4)(MULT_SIZE-1) & MULT_16_3(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(3,4)(MULT_SIZE-1) & MULT_16_4(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(3,4)<=signed(MULT_16_5(3,4)(MULT_SIZE-1) & MULT_16_5(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(3,4)(MULT_SIZE-1) & MULT_16_6(3,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(3,4) ------------------

			MULTS_1_1_1(4,0)<=signed(MULT_1_1(4,0)(MULT_SIZE-1) & MULT_1_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(4,0)(MULT_SIZE-1) & MULT_1_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(4,0)<=signed(MULT_1_3(4,0)(MULT_SIZE-1) & MULT_1_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(4,0)(MULT_SIZE-1) & MULT_1_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(4,0)<=signed(MULT_1_5(4,0)(MULT_SIZE-1) & MULT_1_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(4,0)(MULT_SIZE-1) & MULT_1_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(4,0)<=signed(MULT_2_1(4,0)(MULT_SIZE-1) & MULT_2_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(4,0)(MULT_SIZE-1) & MULT_2_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(4,0)<=signed(MULT_2_3(4,0)(MULT_SIZE-1) & MULT_2_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(4,0)(MULT_SIZE-1) & MULT_2_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(4,0)<=signed(MULT_2_5(4,0)(MULT_SIZE-1) & MULT_2_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(4,0)(MULT_SIZE-1) & MULT_2_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(4,0)<=signed(MULT_3_1(4,0)(MULT_SIZE-1) & MULT_3_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(4,0)(MULT_SIZE-1) & MULT_3_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(4,0)<=signed(MULT_3_3(4,0)(MULT_SIZE-1) & MULT_3_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(4,0)(MULT_SIZE-1) & MULT_3_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(4,0)<=signed(MULT_3_5(4,0)(MULT_SIZE-1) & MULT_3_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(4,0)(MULT_SIZE-1) & MULT_3_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(4,0)<=signed(MULT_4_1(4,0)(MULT_SIZE-1) & MULT_4_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(4,0)(MULT_SIZE-1) & MULT_4_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(4,0)<=signed(MULT_4_3(4,0)(MULT_SIZE-1) & MULT_4_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(4,0)(MULT_SIZE-1) & MULT_4_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(4,0)<=signed(MULT_4_5(4,0)(MULT_SIZE-1) & MULT_4_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(4,0)(MULT_SIZE-1) & MULT_4_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(4,0)<=signed(MULT_5_1(4,0)(MULT_SIZE-1) & MULT_5_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(4,0)(MULT_SIZE-1) & MULT_5_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(4,0)<=signed(MULT_5_3(4,0)(MULT_SIZE-1) & MULT_5_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(4,0)(MULT_SIZE-1) & MULT_5_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(4,0)<=signed(MULT_5_5(4,0)(MULT_SIZE-1) & MULT_5_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(4,0)(MULT_SIZE-1) & MULT_5_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(4,0)<=signed(MULT_6_1(4,0)(MULT_SIZE-1) & MULT_6_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(4,0)(MULT_SIZE-1) & MULT_6_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(4,0)<=signed(MULT_6_3(4,0)(MULT_SIZE-1) & MULT_6_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(4,0)(MULT_SIZE-1) & MULT_6_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(4,0)<=signed(MULT_6_5(4,0)(MULT_SIZE-1) & MULT_6_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(4,0)(MULT_SIZE-1) & MULT_6_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(4,0)<=signed(MULT_7_1(4,0)(MULT_SIZE-1) & MULT_7_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(4,0)(MULT_SIZE-1) & MULT_7_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(4,0)<=signed(MULT_7_3(4,0)(MULT_SIZE-1) & MULT_7_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(4,0)(MULT_SIZE-1) & MULT_7_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(4,0)<=signed(MULT_7_5(4,0)(MULT_SIZE-1) & MULT_7_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(4,0)(MULT_SIZE-1) & MULT_7_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(4,0)<=signed(MULT_8_1(4,0)(MULT_SIZE-1) & MULT_8_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(4,0)(MULT_SIZE-1) & MULT_8_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(4,0)<=signed(MULT_8_3(4,0)(MULT_SIZE-1) & MULT_8_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(4,0)(MULT_SIZE-1) & MULT_8_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(4,0)<=signed(MULT_8_5(4,0)(MULT_SIZE-1) & MULT_8_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(4,0)(MULT_SIZE-1) & MULT_8_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(4,0)<=signed(MULT_9_1(4,0)(MULT_SIZE-1) & MULT_9_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(4,0)(MULT_SIZE-1) & MULT_9_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(4,0)<=signed(MULT_9_3(4,0)(MULT_SIZE-1) & MULT_9_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(4,0)(MULT_SIZE-1) & MULT_9_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(4,0)<=signed(MULT_9_5(4,0)(MULT_SIZE-1) & MULT_9_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(4,0)(MULT_SIZE-1) & MULT_9_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(4,0)<=signed(MULT_10_1(4,0)(MULT_SIZE-1) & MULT_10_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(4,0)(MULT_SIZE-1) & MULT_10_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(4,0)<=signed(MULT_10_3(4,0)(MULT_SIZE-1) & MULT_10_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(4,0)(MULT_SIZE-1) & MULT_10_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(4,0)<=signed(MULT_10_5(4,0)(MULT_SIZE-1) & MULT_10_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(4,0)(MULT_SIZE-1) & MULT_10_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(4,0)<=signed(MULT_11_1(4,0)(MULT_SIZE-1) & MULT_11_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(4,0)(MULT_SIZE-1) & MULT_11_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(4,0)<=signed(MULT_11_3(4,0)(MULT_SIZE-1) & MULT_11_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(4,0)(MULT_SIZE-1) & MULT_11_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(4,0)<=signed(MULT_11_5(4,0)(MULT_SIZE-1) & MULT_11_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(4,0)(MULT_SIZE-1) & MULT_11_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(4,0)<=signed(MULT_12_1(4,0)(MULT_SIZE-1) & MULT_12_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(4,0)(MULT_SIZE-1) & MULT_12_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(4,0)<=signed(MULT_12_3(4,0)(MULT_SIZE-1) & MULT_12_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(4,0)(MULT_SIZE-1) & MULT_12_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(4,0)<=signed(MULT_12_5(4,0)(MULT_SIZE-1) & MULT_12_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(4,0)(MULT_SIZE-1) & MULT_12_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(4,0)<=signed(MULT_13_1(4,0)(MULT_SIZE-1) & MULT_13_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(4,0)(MULT_SIZE-1) & MULT_13_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(4,0)<=signed(MULT_13_3(4,0)(MULT_SIZE-1) & MULT_13_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(4,0)(MULT_SIZE-1) & MULT_13_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(4,0)<=signed(MULT_13_5(4,0)(MULT_SIZE-1) & MULT_13_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(4,0)(MULT_SIZE-1) & MULT_13_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(4,0)<=signed(MULT_14_1(4,0)(MULT_SIZE-1) & MULT_14_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(4,0)(MULT_SIZE-1) & MULT_14_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(4,0)<=signed(MULT_14_3(4,0)(MULT_SIZE-1) & MULT_14_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(4,0)(MULT_SIZE-1) & MULT_14_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(4,0)<=signed(MULT_14_5(4,0)(MULT_SIZE-1) & MULT_14_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(4,0)(MULT_SIZE-1) & MULT_14_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(4,0)<=signed(MULT_15_1(4,0)(MULT_SIZE-1) & MULT_15_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(4,0)(MULT_SIZE-1) & MULT_15_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(4,0)<=signed(MULT_15_3(4,0)(MULT_SIZE-1) & MULT_15_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(4,0)(MULT_SIZE-1) & MULT_15_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(4,0)<=signed(MULT_15_5(4,0)(MULT_SIZE-1) & MULT_15_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(4,0)(MULT_SIZE-1) & MULT_15_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(4,0)<=signed(MULT_16_1(4,0)(MULT_SIZE-1) & MULT_16_1(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(4,0)(MULT_SIZE-1) & MULT_16_2(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(4,0)<=signed(MULT_16_3(4,0)(MULT_SIZE-1) & MULT_16_3(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(4,0)(MULT_SIZE-1) & MULT_16_4(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(4,0)<=signed(MULT_16_5(4,0)(MULT_SIZE-1) & MULT_16_5(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(4,0)(MULT_SIZE-1) & MULT_16_6(4,0)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(4,0) ------------------

			MULTS_1_1_1(4,1)<=signed(MULT_1_1(4,1)(MULT_SIZE-1) & MULT_1_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(4,1)(MULT_SIZE-1) & MULT_1_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(4,1)<=signed(MULT_1_3(4,1)(MULT_SIZE-1) & MULT_1_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(4,1)(MULT_SIZE-1) & MULT_1_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(4,1)<=signed(MULT_1_5(4,1)(MULT_SIZE-1) & MULT_1_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(4,1)(MULT_SIZE-1) & MULT_1_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(4,1)<=signed(MULT_2_1(4,1)(MULT_SIZE-1) & MULT_2_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(4,1)(MULT_SIZE-1) & MULT_2_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(4,1)<=signed(MULT_2_3(4,1)(MULT_SIZE-1) & MULT_2_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(4,1)(MULT_SIZE-1) & MULT_2_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(4,1)<=signed(MULT_2_5(4,1)(MULT_SIZE-1) & MULT_2_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(4,1)(MULT_SIZE-1) & MULT_2_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(4,1)<=signed(MULT_3_1(4,1)(MULT_SIZE-1) & MULT_3_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(4,1)(MULT_SIZE-1) & MULT_3_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(4,1)<=signed(MULT_3_3(4,1)(MULT_SIZE-1) & MULT_3_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(4,1)(MULT_SIZE-1) & MULT_3_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(4,1)<=signed(MULT_3_5(4,1)(MULT_SIZE-1) & MULT_3_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(4,1)(MULT_SIZE-1) & MULT_3_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(4,1)<=signed(MULT_4_1(4,1)(MULT_SIZE-1) & MULT_4_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(4,1)(MULT_SIZE-1) & MULT_4_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(4,1)<=signed(MULT_4_3(4,1)(MULT_SIZE-1) & MULT_4_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(4,1)(MULT_SIZE-1) & MULT_4_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(4,1)<=signed(MULT_4_5(4,1)(MULT_SIZE-1) & MULT_4_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(4,1)(MULT_SIZE-1) & MULT_4_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(4,1)<=signed(MULT_5_1(4,1)(MULT_SIZE-1) & MULT_5_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(4,1)(MULT_SIZE-1) & MULT_5_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(4,1)<=signed(MULT_5_3(4,1)(MULT_SIZE-1) & MULT_5_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(4,1)(MULT_SIZE-1) & MULT_5_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(4,1)<=signed(MULT_5_5(4,1)(MULT_SIZE-1) & MULT_5_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(4,1)(MULT_SIZE-1) & MULT_5_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(4,1)<=signed(MULT_6_1(4,1)(MULT_SIZE-1) & MULT_6_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(4,1)(MULT_SIZE-1) & MULT_6_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(4,1)<=signed(MULT_6_3(4,1)(MULT_SIZE-1) & MULT_6_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(4,1)(MULT_SIZE-1) & MULT_6_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(4,1)<=signed(MULT_6_5(4,1)(MULT_SIZE-1) & MULT_6_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(4,1)(MULT_SIZE-1) & MULT_6_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(4,1)<=signed(MULT_7_1(4,1)(MULT_SIZE-1) & MULT_7_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(4,1)(MULT_SIZE-1) & MULT_7_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(4,1)<=signed(MULT_7_3(4,1)(MULT_SIZE-1) & MULT_7_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(4,1)(MULT_SIZE-1) & MULT_7_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(4,1)<=signed(MULT_7_5(4,1)(MULT_SIZE-1) & MULT_7_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(4,1)(MULT_SIZE-1) & MULT_7_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(4,1)<=signed(MULT_8_1(4,1)(MULT_SIZE-1) & MULT_8_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(4,1)(MULT_SIZE-1) & MULT_8_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(4,1)<=signed(MULT_8_3(4,1)(MULT_SIZE-1) & MULT_8_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(4,1)(MULT_SIZE-1) & MULT_8_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(4,1)<=signed(MULT_8_5(4,1)(MULT_SIZE-1) & MULT_8_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(4,1)(MULT_SIZE-1) & MULT_8_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(4,1)<=signed(MULT_9_1(4,1)(MULT_SIZE-1) & MULT_9_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(4,1)(MULT_SIZE-1) & MULT_9_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(4,1)<=signed(MULT_9_3(4,1)(MULT_SIZE-1) & MULT_9_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(4,1)(MULT_SIZE-1) & MULT_9_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(4,1)<=signed(MULT_9_5(4,1)(MULT_SIZE-1) & MULT_9_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(4,1)(MULT_SIZE-1) & MULT_9_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(4,1)<=signed(MULT_10_1(4,1)(MULT_SIZE-1) & MULT_10_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(4,1)(MULT_SIZE-1) & MULT_10_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(4,1)<=signed(MULT_10_3(4,1)(MULT_SIZE-1) & MULT_10_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(4,1)(MULT_SIZE-1) & MULT_10_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(4,1)<=signed(MULT_10_5(4,1)(MULT_SIZE-1) & MULT_10_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(4,1)(MULT_SIZE-1) & MULT_10_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(4,1)<=signed(MULT_11_1(4,1)(MULT_SIZE-1) & MULT_11_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(4,1)(MULT_SIZE-1) & MULT_11_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(4,1)<=signed(MULT_11_3(4,1)(MULT_SIZE-1) & MULT_11_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(4,1)(MULT_SIZE-1) & MULT_11_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(4,1)<=signed(MULT_11_5(4,1)(MULT_SIZE-1) & MULT_11_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(4,1)(MULT_SIZE-1) & MULT_11_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(4,1)<=signed(MULT_12_1(4,1)(MULT_SIZE-1) & MULT_12_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(4,1)(MULT_SIZE-1) & MULT_12_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(4,1)<=signed(MULT_12_3(4,1)(MULT_SIZE-1) & MULT_12_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(4,1)(MULT_SIZE-1) & MULT_12_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(4,1)<=signed(MULT_12_5(4,1)(MULT_SIZE-1) & MULT_12_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(4,1)(MULT_SIZE-1) & MULT_12_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(4,1)<=signed(MULT_13_1(4,1)(MULT_SIZE-1) & MULT_13_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(4,1)(MULT_SIZE-1) & MULT_13_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(4,1)<=signed(MULT_13_3(4,1)(MULT_SIZE-1) & MULT_13_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(4,1)(MULT_SIZE-1) & MULT_13_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(4,1)<=signed(MULT_13_5(4,1)(MULT_SIZE-1) & MULT_13_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(4,1)(MULT_SIZE-1) & MULT_13_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(4,1)<=signed(MULT_14_1(4,1)(MULT_SIZE-1) & MULT_14_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(4,1)(MULT_SIZE-1) & MULT_14_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(4,1)<=signed(MULT_14_3(4,1)(MULT_SIZE-1) & MULT_14_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(4,1)(MULT_SIZE-1) & MULT_14_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(4,1)<=signed(MULT_14_5(4,1)(MULT_SIZE-1) & MULT_14_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(4,1)(MULT_SIZE-1) & MULT_14_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(4,1)<=signed(MULT_15_1(4,1)(MULT_SIZE-1) & MULT_15_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(4,1)(MULT_SIZE-1) & MULT_15_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(4,1)<=signed(MULT_15_3(4,1)(MULT_SIZE-1) & MULT_15_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(4,1)(MULT_SIZE-1) & MULT_15_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(4,1)<=signed(MULT_15_5(4,1)(MULT_SIZE-1) & MULT_15_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(4,1)(MULT_SIZE-1) & MULT_15_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(4,1)<=signed(MULT_16_1(4,1)(MULT_SIZE-1) & MULT_16_1(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(4,1)(MULT_SIZE-1) & MULT_16_2(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(4,1)<=signed(MULT_16_3(4,1)(MULT_SIZE-1) & MULT_16_3(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(4,1)(MULT_SIZE-1) & MULT_16_4(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(4,1)<=signed(MULT_16_5(4,1)(MULT_SIZE-1) & MULT_16_5(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(4,1)(MULT_SIZE-1) & MULT_16_6(4,1)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(4,1) ------------------

			MULTS_1_1_1(4,2)<=signed(MULT_1_1(4,2)(MULT_SIZE-1) & MULT_1_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(4,2)(MULT_SIZE-1) & MULT_1_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(4,2)<=signed(MULT_1_3(4,2)(MULT_SIZE-1) & MULT_1_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(4,2)(MULT_SIZE-1) & MULT_1_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(4,2)<=signed(MULT_1_5(4,2)(MULT_SIZE-1) & MULT_1_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(4,2)(MULT_SIZE-1) & MULT_1_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(4,2)<=signed(MULT_2_1(4,2)(MULT_SIZE-1) & MULT_2_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(4,2)(MULT_SIZE-1) & MULT_2_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(4,2)<=signed(MULT_2_3(4,2)(MULT_SIZE-1) & MULT_2_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(4,2)(MULT_SIZE-1) & MULT_2_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(4,2)<=signed(MULT_2_5(4,2)(MULT_SIZE-1) & MULT_2_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(4,2)(MULT_SIZE-1) & MULT_2_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(4,2)<=signed(MULT_3_1(4,2)(MULT_SIZE-1) & MULT_3_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(4,2)(MULT_SIZE-1) & MULT_3_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(4,2)<=signed(MULT_3_3(4,2)(MULT_SIZE-1) & MULT_3_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(4,2)(MULT_SIZE-1) & MULT_3_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(4,2)<=signed(MULT_3_5(4,2)(MULT_SIZE-1) & MULT_3_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(4,2)(MULT_SIZE-1) & MULT_3_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(4,2)<=signed(MULT_4_1(4,2)(MULT_SIZE-1) & MULT_4_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(4,2)(MULT_SIZE-1) & MULT_4_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(4,2)<=signed(MULT_4_3(4,2)(MULT_SIZE-1) & MULT_4_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(4,2)(MULT_SIZE-1) & MULT_4_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(4,2)<=signed(MULT_4_5(4,2)(MULT_SIZE-1) & MULT_4_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(4,2)(MULT_SIZE-1) & MULT_4_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(4,2)<=signed(MULT_5_1(4,2)(MULT_SIZE-1) & MULT_5_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(4,2)(MULT_SIZE-1) & MULT_5_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(4,2)<=signed(MULT_5_3(4,2)(MULT_SIZE-1) & MULT_5_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(4,2)(MULT_SIZE-1) & MULT_5_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(4,2)<=signed(MULT_5_5(4,2)(MULT_SIZE-1) & MULT_5_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(4,2)(MULT_SIZE-1) & MULT_5_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(4,2)<=signed(MULT_6_1(4,2)(MULT_SIZE-1) & MULT_6_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(4,2)(MULT_SIZE-1) & MULT_6_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(4,2)<=signed(MULT_6_3(4,2)(MULT_SIZE-1) & MULT_6_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(4,2)(MULT_SIZE-1) & MULT_6_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(4,2)<=signed(MULT_6_5(4,2)(MULT_SIZE-1) & MULT_6_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(4,2)(MULT_SIZE-1) & MULT_6_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(4,2)<=signed(MULT_7_1(4,2)(MULT_SIZE-1) & MULT_7_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(4,2)(MULT_SIZE-1) & MULT_7_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(4,2)<=signed(MULT_7_3(4,2)(MULT_SIZE-1) & MULT_7_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(4,2)(MULT_SIZE-1) & MULT_7_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(4,2)<=signed(MULT_7_5(4,2)(MULT_SIZE-1) & MULT_7_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(4,2)(MULT_SIZE-1) & MULT_7_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(4,2)<=signed(MULT_8_1(4,2)(MULT_SIZE-1) & MULT_8_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(4,2)(MULT_SIZE-1) & MULT_8_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(4,2)<=signed(MULT_8_3(4,2)(MULT_SIZE-1) & MULT_8_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(4,2)(MULT_SIZE-1) & MULT_8_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(4,2)<=signed(MULT_8_5(4,2)(MULT_SIZE-1) & MULT_8_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(4,2)(MULT_SIZE-1) & MULT_8_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(4,2)<=signed(MULT_9_1(4,2)(MULT_SIZE-1) & MULT_9_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(4,2)(MULT_SIZE-1) & MULT_9_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(4,2)<=signed(MULT_9_3(4,2)(MULT_SIZE-1) & MULT_9_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(4,2)(MULT_SIZE-1) & MULT_9_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(4,2)<=signed(MULT_9_5(4,2)(MULT_SIZE-1) & MULT_9_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(4,2)(MULT_SIZE-1) & MULT_9_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(4,2)<=signed(MULT_10_1(4,2)(MULT_SIZE-1) & MULT_10_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(4,2)(MULT_SIZE-1) & MULT_10_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(4,2)<=signed(MULT_10_3(4,2)(MULT_SIZE-1) & MULT_10_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(4,2)(MULT_SIZE-1) & MULT_10_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(4,2)<=signed(MULT_10_5(4,2)(MULT_SIZE-1) & MULT_10_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(4,2)(MULT_SIZE-1) & MULT_10_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(4,2)<=signed(MULT_11_1(4,2)(MULT_SIZE-1) & MULT_11_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(4,2)(MULT_SIZE-1) & MULT_11_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(4,2)<=signed(MULT_11_3(4,2)(MULT_SIZE-1) & MULT_11_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(4,2)(MULT_SIZE-1) & MULT_11_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(4,2)<=signed(MULT_11_5(4,2)(MULT_SIZE-1) & MULT_11_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(4,2)(MULT_SIZE-1) & MULT_11_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(4,2)<=signed(MULT_12_1(4,2)(MULT_SIZE-1) & MULT_12_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(4,2)(MULT_SIZE-1) & MULT_12_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(4,2)<=signed(MULT_12_3(4,2)(MULT_SIZE-1) & MULT_12_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(4,2)(MULT_SIZE-1) & MULT_12_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(4,2)<=signed(MULT_12_5(4,2)(MULT_SIZE-1) & MULT_12_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(4,2)(MULT_SIZE-1) & MULT_12_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(4,2)<=signed(MULT_13_1(4,2)(MULT_SIZE-1) & MULT_13_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(4,2)(MULT_SIZE-1) & MULT_13_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(4,2)<=signed(MULT_13_3(4,2)(MULT_SIZE-1) & MULT_13_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(4,2)(MULT_SIZE-1) & MULT_13_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(4,2)<=signed(MULT_13_5(4,2)(MULT_SIZE-1) & MULT_13_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(4,2)(MULT_SIZE-1) & MULT_13_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(4,2)<=signed(MULT_14_1(4,2)(MULT_SIZE-1) & MULT_14_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(4,2)(MULT_SIZE-1) & MULT_14_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(4,2)<=signed(MULT_14_3(4,2)(MULT_SIZE-1) & MULT_14_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(4,2)(MULT_SIZE-1) & MULT_14_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(4,2)<=signed(MULT_14_5(4,2)(MULT_SIZE-1) & MULT_14_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(4,2)(MULT_SIZE-1) & MULT_14_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(4,2)<=signed(MULT_15_1(4,2)(MULT_SIZE-1) & MULT_15_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(4,2)(MULT_SIZE-1) & MULT_15_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(4,2)<=signed(MULT_15_3(4,2)(MULT_SIZE-1) & MULT_15_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(4,2)(MULT_SIZE-1) & MULT_15_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(4,2)<=signed(MULT_15_5(4,2)(MULT_SIZE-1) & MULT_15_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(4,2)(MULT_SIZE-1) & MULT_15_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(4,2)<=signed(MULT_16_1(4,2)(MULT_SIZE-1) & MULT_16_1(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(4,2)(MULT_SIZE-1) & MULT_16_2(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(4,2)<=signed(MULT_16_3(4,2)(MULT_SIZE-1) & MULT_16_3(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(4,2)(MULT_SIZE-1) & MULT_16_4(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(4,2)<=signed(MULT_16_5(4,2)(MULT_SIZE-1) & MULT_16_5(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(4,2)(MULT_SIZE-1) & MULT_16_6(4,2)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(4,2) ------------------

			MULTS_1_1_1(4,3)<=signed(MULT_1_1(4,3)(MULT_SIZE-1) & MULT_1_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(4,3)(MULT_SIZE-1) & MULT_1_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(4,3)<=signed(MULT_1_3(4,3)(MULT_SIZE-1) & MULT_1_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(4,3)(MULT_SIZE-1) & MULT_1_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(4,3)<=signed(MULT_1_5(4,3)(MULT_SIZE-1) & MULT_1_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(4,3)(MULT_SIZE-1) & MULT_1_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(4,3)<=signed(MULT_2_1(4,3)(MULT_SIZE-1) & MULT_2_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(4,3)(MULT_SIZE-1) & MULT_2_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(4,3)<=signed(MULT_2_3(4,3)(MULT_SIZE-1) & MULT_2_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(4,3)(MULT_SIZE-1) & MULT_2_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(4,3)<=signed(MULT_2_5(4,3)(MULT_SIZE-1) & MULT_2_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(4,3)(MULT_SIZE-1) & MULT_2_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(4,3)<=signed(MULT_3_1(4,3)(MULT_SIZE-1) & MULT_3_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(4,3)(MULT_SIZE-1) & MULT_3_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(4,3)<=signed(MULT_3_3(4,3)(MULT_SIZE-1) & MULT_3_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(4,3)(MULT_SIZE-1) & MULT_3_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(4,3)<=signed(MULT_3_5(4,3)(MULT_SIZE-1) & MULT_3_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(4,3)(MULT_SIZE-1) & MULT_3_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(4,3)<=signed(MULT_4_1(4,3)(MULT_SIZE-1) & MULT_4_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(4,3)(MULT_SIZE-1) & MULT_4_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(4,3)<=signed(MULT_4_3(4,3)(MULT_SIZE-1) & MULT_4_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(4,3)(MULT_SIZE-1) & MULT_4_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(4,3)<=signed(MULT_4_5(4,3)(MULT_SIZE-1) & MULT_4_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(4,3)(MULT_SIZE-1) & MULT_4_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(4,3)<=signed(MULT_5_1(4,3)(MULT_SIZE-1) & MULT_5_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(4,3)(MULT_SIZE-1) & MULT_5_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(4,3)<=signed(MULT_5_3(4,3)(MULT_SIZE-1) & MULT_5_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(4,3)(MULT_SIZE-1) & MULT_5_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(4,3)<=signed(MULT_5_5(4,3)(MULT_SIZE-1) & MULT_5_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(4,3)(MULT_SIZE-1) & MULT_5_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(4,3)<=signed(MULT_6_1(4,3)(MULT_SIZE-1) & MULT_6_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(4,3)(MULT_SIZE-1) & MULT_6_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(4,3)<=signed(MULT_6_3(4,3)(MULT_SIZE-1) & MULT_6_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(4,3)(MULT_SIZE-1) & MULT_6_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(4,3)<=signed(MULT_6_5(4,3)(MULT_SIZE-1) & MULT_6_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(4,3)(MULT_SIZE-1) & MULT_6_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(4,3)<=signed(MULT_7_1(4,3)(MULT_SIZE-1) & MULT_7_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(4,3)(MULT_SIZE-1) & MULT_7_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(4,3)<=signed(MULT_7_3(4,3)(MULT_SIZE-1) & MULT_7_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(4,3)(MULT_SIZE-1) & MULT_7_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(4,3)<=signed(MULT_7_5(4,3)(MULT_SIZE-1) & MULT_7_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(4,3)(MULT_SIZE-1) & MULT_7_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(4,3)<=signed(MULT_8_1(4,3)(MULT_SIZE-1) & MULT_8_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(4,3)(MULT_SIZE-1) & MULT_8_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(4,3)<=signed(MULT_8_3(4,3)(MULT_SIZE-1) & MULT_8_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(4,3)(MULT_SIZE-1) & MULT_8_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(4,3)<=signed(MULT_8_5(4,3)(MULT_SIZE-1) & MULT_8_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(4,3)(MULT_SIZE-1) & MULT_8_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(4,3)<=signed(MULT_9_1(4,3)(MULT_SIZE-1) & MULT_9_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(4,3)(MULT_SIZE-1) & MULT_9_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(4,3)<=signed(MULT_9_3(4,3)(MULT_SIZE-1) & MULT_9_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(4,3)(MULT_SIZE-1) & MULT_9_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(4,3)<=signed(MULT_9_5(4,3)(MULT_SIZE-1) & MULT_9_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(4,3)(MULT_SIZE-1) & MULT_9_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(4,3)<=signed(MULT_10_1(4,3)(MULT_SIZE-1) & MULT_10_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(4,3)(MULT_SIZE-1) & MULT_10_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(4,3)<=signed(MULT_10_3(4,3)(MULT_SIZE-1) & MULT_10_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(4,3)(MULT_SIZE-1) & MULT_10_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(4,3)<=signed(MULT_10_5(4,3)(MULT_SIZE-1) & MULT_10_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(4,3)(MULT_SIZE-1) & MULT_10_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(4,3)<=signed(MULT_11_1(4,3)(MULT_SIZE-1) & MULT_11_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(4,3)(MULT_SIZE-1) & MULT_11_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(4,3)<=signed(MULT_11_3(4,3)(MULT_SIZE-1) & MULT_11_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(4,3)(MULT_SIZE-1) & MULT_11_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(4,3)<=signed(MULT_11_5(4,3)(MULT_SIZE-1) & MULT_11_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(4,3)(MULT_SIZE-1) & MULT_11_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(4,3)<=signed(MULT_12_1(4,3)(MULT_SIZE-1) & MULT_12_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(4,3)(MULT_SIZE-1) & MULT_12_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(4,3)<=signed(MULT_12_3(4,3)(MULT_SIZE-1) & MULT_12_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(4,3)(MULT_SIZE-1) & MULT_12_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(4,3)<=signed(MULT_12_5(4,3)(MULT_SIZE-1) & MULT_12_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(4,3)(MULT_SIZE-1) & MULT_12_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(4,3)<=signed(MULT_13_1(4,3)(MULT_SIZE-1) & MULT_13_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(4,3)(MULT_SIZE-1) & MULT_13_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(4,3)<=signed(MULT_13_3(4,3)(MULT_SIZE-1) & MULT_13_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(4,3)(MULT_SIZE-1) & MULT_13_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(4,3)<=signed(MULT_13_5(4,3)(MULT_SIZE-1) & MULT_13_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(4,3)(MULT_SIZE-1) & MULT_13_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(4,3)<=signed(MULT_14_1(4,3)(MULT_SIZE-1) & MULT_14_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(4,3)(MULT_SIZE-1) & MULT_14_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(4,3)<=signed(MULT_14_3(4,3)(MULT_SIZE-1) & MULT_14_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(4,3)(MULT_SIZE-1) & MULT_14_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(4,3)<=signed(MULT_14_5(4,3)(MULT_SIZE-1) & MULT_14_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(4,3)(MULT_SIZE-1) & MULT_14_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(4,3)<=signed(MULT_15_1(4,3)(MULT_SIZE-1) & MULT_15_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(4,3)(MULT_SIZE-1) & MULT_15_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(4,3)<=signed(MULT_15_3(4,3)(MULT_SIZE-1) & MULT_15_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(4,3)(MULT_SIZE-1) & MULT_15_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(4,3)<=signed(MULT_15_5(4,3)(MULT_SIZE-1) & MULT_15_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(4,3)(MULT_SIZE-1) & MULT_15_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(4,3)<=signed(MULT_16_1(4,3)(MULT_SIZE-1) & MULT_16_1(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(4,3)(MULT_SIZE-1) & MULT_16_2(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(4,3)<=signed(MULT_16_3(4,3)(MULT_SIZE-1) & MULT_16_3(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(4,3)(MULT_SIZE-1) & MULT_16_4(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(4,3)<=signed(MULT_16_5(4,3)(MULT_SIZE-1) & MULT_16_5(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(4,3)(MULT_SIZE-1) & MULT_16_6(4,3)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(4,3) ------------------

			MULTS_1_1_1(4,4)<=signed(MULT_1_1(4,4)(MULT_SIZE-1) & MULT_1_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_2(4,4)(MULT_SIZE-1) & MULT_1_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_2(4,4)<=signed(MULT_1_3(4,4)(MULT_SIZE-1) & MULT_1_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_4(4,4)(MULT_SIZE-1) & MULT_1_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_1_3(4,4)<=signed(MULT_1_5(4,4)(MULT_SIZE-1) & MULT_1_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_1_6(4,4)(MULT_SIZE-1) & MULT_1_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_1_2_1(4,4)<=signed(MULT_2_1(4,4)(MULT_SIZE-1) & MULT_2_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_2(4,4)(MULT_SIZE-1) & MULT_2_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_2(4,4)<=signed(MULT_2_3(4,4)(MULT_SIZE-1) & MULT_2_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_4(4,4)(MULT_SIZE-1) & MULT_2_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_2_3(4,4)<=signed(MULT_2_5(4,4)(MULT_SIZE-1) & MULT_2_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_2_6(4,4)(MULT_SIZE-1) & MULT_2_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_1_3_1(4,4)<=signed(MULT_3_1(4,4)(MULT_SIZE-1) & MULT_3_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_2(4,4)(MULT_SIZE-1) & MULT_3_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_2(4,4)<=signed(MULT_3_3(4,4)(MULT_SIZE-1) & MULT_3_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_4(4,4)(MULT_SIZE-1) & MULT_3_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_3_3(4,4)<=signed(MULT_3_5(4,4)(MULT_SIZE-1) & MULT_3_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_3_6(4,4)(MULT_SIZE-1) & MULT_3_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_1_4_1(4,4)<=signed(MULT_4_1(4,4)(MULT_SIZE-1) & MULT_4_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_2(4,4)(MULT_SIZE-1) & MULT_4_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_2(4,4)<=signed(MULT_4_3(4,4)(MULT_SIZE-1) & MULT_4_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_4(4,4)(MULT_SIZE-1) & MULT_4_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_4_3(4,4)<=signed(MULT_4_5(4,4)(MULT_SIZE-1) & MULT_4_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_4_6(4,4)(MULT_SIZE-1) & MULT_4_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_1_5_1(4,4)<=signed(MULT_5_1(4,4)(MULT_SIZE-1) & MULT_5_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_2(4,4)(MULT_SIZE-1) & MULT_5_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_2(4,4)<=signed(MULT_5_3(4,4)(MULT_SIZE-1) & MULT_5_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_4(4,4)(MULT_SIZE-1) & MULT_5_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_5_3(4,4)<=signed(MULT_5_5(4,4)(MULT_SIZE-1) & MULT_5_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_5_6(4,4)(MULT_SIZE-1) & MULT_5_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_1_6_1(4,4)<=signed(MULT_6_1(4,4)(MULT_SIZE-1) & MULT_6_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_2(4,4)(MULT_SIZE-1) & MULT_6_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_2(4,4)<=signed(MULT_6_3(4,4)(MULT_SIZE-1) & MULT_6_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_4(4,4)(MULT_SIZE-1) & MULT_6_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_6_3(4,4)<=signed(MULT_6_5(4,4)(MULT_SIZE-1) & MULT_6_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_6_6(4,4)(MULT_SIZE-1) & MULT_6_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_1_7_1(4,4)<=signed(MULT_7_1(4,4)(MULT_SIZE-1) & MULT_7_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_2(4,4)(MULT_SIZE-1) & MULT_7_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_2(4,4)<=signed(MULT_7_3(4,4)(MULT_SIZE-1) & MULT_7_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_4(4,4)(MULT_SIZE-1) & MULT_7_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_7_3(4,4)<=signed(MULT_7_5(4,4)(MULT_SIZE-1) & MULT_7_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_7_6(4,4)(MULT_SIZE-1) & MULT_7_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_1_8_1(4,4)<=signed(MULT_8_1(4,4)(MULT_SIZE-1) & MULT_8_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_2(4,4)(MULT_SIZE-1) & MULT_8_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_2(4,4)<=signed(MULT_8_3(4,4)(MULT_SIZE-1) & MULT_8_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_4(4,4)(MULT_SIZE-1) & MULT_8_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_8_3(4,4)<=signed(MULT_8_5(4,4)(MULT_SIZE-1) & MULT_8_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_8_6(4,4)(MULT_SIZE-1) & MULT_8_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_1_9_1(4,4)<=signed(MULT_9_1(4,4)(MULT_SIZE-1) & MULT_9_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_2(4,4)(MULT_SIZE-1) & MULT_9_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_2(4,4)<=signed(MULT_9_3(4,4)(MULT_SIZE-1) & MULT_9_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_4(4,4)(MULT_SIZE-1) & MULT_9_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_9_3(4,4)<=signed(MULT_9_5(4,4)(MULT_SIZE-1) & MULT_9_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_9_6(4,4)(MULT_SIZE-1) & MULT_9_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_1_10_1(4,4)<=signed(MULT_10_1(4,4)(MULT_SIZE-1) & MULT_10_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_2(4,4)(MULT_SIZE-1) & MULT_10_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_2(4,4)<=signed(MULT_10_3(4,4)(MULT_SIZE-1) & MULT_10_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_4(4,4)(MULT_SIZE-1) & MULT_10_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_10_3(4,4)<=signed(MULT_10_5(4,4)(MULT_SIZE-1) & MULT_10_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_10_6(4,4)(MULT_SIZE-1) & MULT_10_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_1_11_1(4,4)<=signed(MULT_11_1(4,4)(MULT_SIZE-1) & MULT_11_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_2(4,4)(MULT_SIZE-1) & MULT_11_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_2(4,4)<=signed(MULT_11_3(4,4)(MULT_SIZE-1) & MULT_11_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_4(4,4)(MULT_SIZE-1) & MULT_11_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_11_3(4,4)<=signed(MULT_11_5(4,4)(MULT_SIZE-1) & MULT_11_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_11_6(4,4)(MULT_SIZE-1) & MULT_11_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_1_12_1(4,4)<=signed(MULT_12_1(4,4)(MULT_SIZE-1) & MULT_12_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_2(4,4)(MULT_SIZE-1) & MULT_12_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_2(4,4)<=signed(MULT_12_3(4,4)(MULT_SIZE-1) & MULT_12_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_4(4,4)(MULT_SIZE-1) & MULT_12_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_12_3(4,4)<=signed(MULT_12_5(4,4)(MULT_SIZE-1) & MULT_12_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_12_6(4,4)(MULT_SIZE-1) & MULT_12_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_1_13_1(4,4)<=signed(MULT_13_1(4,4)(MULT_SIZE-1) & MULT_13_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_2(4,4)(MULT_SIZE-1) & MULT_13_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_2(4,4)<=signed(MULT_13_3(4,4)(MULT_SIZE-1) & MULT_13_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_4(4,4)(MULT_SIZE-1) & MULT_13_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_13_3(4,4)<=signed(MULT_13_5(4,4)(MULT_SIZE-1) & MULT_13_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_13_6(4,4)(MULT_SIZE-1) & MULT_13_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_1_14_1(4,4)<=signed(MULT_14_1(4,4)(MULT_SIZE-1) & MULT_14_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_2(4,4)(MULT_SIZE-1) & MULT_14_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_2(4,4)<=signed(MULT_14_3(4,4)(MULT_SIZE-1) & MULT_14_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_4(4,4)(MULT_SIZE-1) & MULT_14_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_14_3(4,4)<=signed(MULT_14_5(4,4)(MULT_SIZE-1) & MULT_14_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_14_6(4,4)(MULT_SIZE-1) & MULT_14_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_1_15_1(4,4)<=signed(MULT_15_1(4,4)(MULT_SIZE-1) & MULT_15_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_2(4,4)(MULT_SIZE-1) & MULT_15_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_2(4,4)<=signed(MULT_15_3(4,4)(MULT_SIZE-1) & MULT_15_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_4(4,4)(MULT_SIZE-1) & MULT_15_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_15_3(4,4)<=signed(MULT_15_5(4,4)(MULT_SIZE-1) & MULT_15_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_15_6(4,4)(MULT_SIZE-1) & MULT_15_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_1_16_1(4,4)<=signed(MULT_16_1(4,4)(MULT_SIZE-1) & MULT_16_1(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_2(4,4)(MULT_SIZE-1) & MULT_16_2(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_2(4,4)<=signed(MULT_16_3(4,4)(MULT_SIZE-1) & MULT_16_3(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_4(4,4)(MULT_SIZE-1) & MULT_16_4(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			MULTS_1_16_3(4,4)<=signed(MULT_16_5(4,4)(MULT_SIZE-1) & MULT_16_5(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2)) + signed(MULT_16_6(4,4)(MULT_SIZE-1) & MULT_16_6(4,4)(MULT_SIZE-3 downto MULT_SIZE-PERCISION-2));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(4,4) ------------------



                     EN_SUM_MULT_2<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_2 = '1' then
			------------------------------------STAGE-2--------------------------------------
			MULTS_2_1_1(0,0)<=signed(MULTS_1_1_1(0,0)(PERCISION) & MULTS_1_1_1(0,0)(PERCISION downto 1));
			MULTS_2_2_1(0,0)<=signed(MULTS_1_2_1(0,0)(PERCISION) & MULTS_1_2_1(0,0)(PERCISION downto 1));
			MULTS_2_3_1(0,0)<=signed(MULTS_1_3_1(0,0)(PERCISION) & MULTS_1_3_1(0,0)(PERCISION downto 1));
			MULTS_2_4_1(0,0)<=signed(MULTS_1_4_1(0,0)(PERCISION) & MULTS_1_4_1(0,0)(PERCISION downto 1));
			MULTS_2_5_1(0,0)<=signed(MULTS_1_5_1(0,0)(PERCISION) & MULTS_1_5_1(0,0)(PERCISION downto 1));
			MULTS_2_6_1(0,0)<=signed(MULTS_1_6_1(0,0)(PERCISION) & MULTS_1_6_1(0,0)(PERCISION downto 1));
			MULTS_2_7_1(0,0)<=signed(MULTS_1_7_1(0,0)(PERCISION) & MULTS_1_7_1(0,0)(PERCISION downto 1));
			MULTS_2_8_1(0,0)<=signed(MULTS_1_8_1(0,0)(PERCISION) & MULTS_1_8_1(0,0)(PERCISION downto 1));
			MULTS_2_9_1(0,0)<=signed(MULTS_1_9_1(0,0)(PERCISION) & MULTS_1_9_1(0,0)(PERCISION downto 1));
			MULTS_2_10_1(0,0)<=signed(MULTS_1_10_1(0,0)(PERCISION) & MULTS_1_10_1(0,0)(PERCISION downto 1));
			MULTS_2_11_1(0,0)<=signed(MULTS_1_11_1(0,0)(PERCISION) & MULTS_1_11_1(0,0)(PERCISION downto 1));
			MULTS_2_12_1(0,0)<=signed(MULTS_1_12_1(0,0)(PERCISION) & MULTS_1_12_1(0,0)(PERCISION downto 1));
			MULTS_2_13_1(0,0)<=signed(MULTS_1_13_1(0,0)(PERCISION) & MULTS_1_13_1(0,0)(PERCISION downto 1));
			MULTS_2_14_1(0,0)<=signed(MULTS_1_14_1(0,0)(PERCISION) & MULTS_1_14_1(0,0)(PERCISION downto 1));
			MULTS_2_15_1(0,0)<=signed(MULTS_1_15_1(0,0)(PERCISION) & MULTS_1_15_1(0,0)(PERCISION downto 1));
			MULTS_2_16_1(0,0)<=signed(MULTS_1_16_1(0,0)(PERCISION) & MULTS_1_16_1(0,0)(PERCISION downto 1));

			MULTS_2_1_1(0,1)<=signed(MULTS_1_1_1(0,1)(PERCISION) & MULTS_1_1_1(0,1)(PERCISION downto 1));
			MULTS_2_2_1(0,1)<=signed(MULTS_1_2_1(0,1)(PERCISION) & MULTS_1_2_1(0,1)(PERCISION downto 1));
			MULTS_2_3_1(0,1)<=signed(MULTS_1_3_1(0,1)(PERCISION) & MULTS_1_3_1(0,1)(PERCISION downto 1));
			MULTS_2_4_1(0,1)<=signed(MULTS_1_4_1(0,1)(PERCISION) & MULTS_1_4_1(0,1)(PERCISION downto 1));
			MULTS_2_5_1(0,1)<=signed(MULTS_1_5_1(0,1)(PERCISION) & MULTS_1_5_1(0,1)(PERCISION downto 1));
			MULTS_2_6_1(0,1)<=signed(MULTS_1_6_1(0,1)(PERCISION) & MULTS_1_6_1(0,1)(PERCISION downto 1));
			MULTS_2_7_1(0,1)<=signed(MULTS_1_7_1(0,1)(PERCISION) & MULTS_1_7_1(0,1)(PERCISION downto 1));
			MULTS_2_8_1(0,1)<=signed(MULTS_1_8_1(0,1)(PERCISION) & MULTS_1_8_1(0,1)(PERCISION downto 1));
			MULTS_2_9_1(0,1)<=signed(MULTS_1_9_1(0,1)(PERCISION) & MULTS_1_9_1(0,1)(PERCISION downto 1));
			MULTS_2_10_1(0,1)<=signed(MULTS_1_10_1(0,1)(PERCISION) & MULTS_1_10_1(0,1)(PERCISION downto 1));
			MULTS_2_11_1(0,1)<=signed(MULTS_1_11_1(0,1)(PERCISION) & MULTS_1_11_1(0,1)(PERCISION downto 1));
			MULTS_2_12_1(0,1)<=signed(MULTS_1_12_1(0,1)(PERCISION) & MULTS_1_12_1(0,1)(PERCISION downto 1));
			MULTS_2_13_1(0,1)<=signed(MULTS_1_13_1(0,1)(PERCISION) & MULTS_1_13_1(0,1)(PERCISION downto 1));
			MULTS_2_14_1(0,1)<=signed(MULTS_1_14_1(0,1)(PERCISION) & MULTS_1_14_1(0,1)(PERCISION downto 1));
			MULTS_2_15_1(0,1)<=signed(MULTS_1_15_1(0,1)(PERCISION) & MULTS_1_15_1(0,1)(PERCISION downto 1));
			MULTS_2_16_1(0,1)<=signed(MULTS_1_16_1(0,1)(PERCISION) & MULTS_1_16_1(0,1)(PERCISION downto 1));

			MULTS_2_1_1(0,2)<=signed(MULTS_1_1_1(0,2)(PERCISION) & MULTS_1_1_1(0,2)(PERCISION downto 1));
			MULTS_2_2_1(0,2)<=signed(MULTS_1_2_1(0,2)(PERCISION) & MULTS_1_2_1(0,2)(PERCISION downto 1));
			MULTS_2_3_1(0,2)<=signed(MULTS_1_3_1(0,2)(PERCISION) & MULTS_1_3_1(0,2)(PERCISION downto 1));
			MULTS_2_4_1(0,2)<=signed(MULTS_1_4_1(0,2)(PERCISION) & MULTS_1_4_1(0,2)(PERCISION downto 1));
			MULTS_2_5_1(0,2)<=signed(MULTS_1_5_1(0,2)(PERCISION) & MULTS_1_5_1(0,2)(PERCISION downto 1));
			MULTS_2_6_1(0,2)<=signed(MULTS_1_6_1(0,2)(PERCISION) & MULTS_1_6_1(0,2)(PERCISION downto 1));
			MULTS_2_7_1(0,2)<=signed(MULTS_1_7_1(0,2)(PERCISION) & MULTS_1_7_1(0,2)(PERCISION downto 1));
			MULTS_2_8_1(0,2)<=signed(MULTS_1_8_1(0,2)(PERCISION) & MULTS_1_8_1(0,2)(PERCISION downto 1));
			MULTS_2_9_1(0,2)<=signed(MULTS_1_9_1(0,2)(PERCISION) & MULTS_1_9_1(0,2)(PERCISION downto 1));
			MULTS_2_10_1(0,2)<=signed(MULTS_1_10_1(0,2)(PERCISION) & MULTS_1_10_1(0,2)(PERCISION downto 1));
			MULTS_2_11_1(0,2)<=signed(MULTS_1_11_1(0,2)(PERCISION) & MULTS_1_11_1(0,2)(PERCISION downto 1));
			MULTS_2_12_1(0,2)<=signed(MULTS_1_12_1(0,2)(PERCISION) & MULTS_1_12_1(0,2)(PERCISION downto 1));
			MULTS_2_13_1(0,2)<=signed(MULTS_1_13_1(0,2)(PERCISION) & MULTS_1_13_1(0,2)(PERCISION downto 1));
			MULTS_2_14_1(0,2)<=signed(MULTS_1_14_1(0,2)(PERCISION) & MULTS_1_14_1(0,2)(PERCISION downto 1));
			MULTS_2_15_1(0,2)<=signed(MULTS_1_15_1(0,2)(PERCISION) & MULTS_1_15_1(0,2)(PERCISION downto 1));
			MULTS_2_16_1(0,2)<=signed(MULTS_1_16_1(0,2)(PERCISION) & MULTS_1_16_1(0,2)(PERCISION downto 1));

			MULTS_2_1_1(0,3)<=signed(MULTS_1_1_1(0,3)(PERCISION) & MULTS_1_1_1(0,3)(PERCISION downto 1));
			MULTS_2_2_1(0,3)<=signed(MULTS_1_2_1(0,3)(PERCISION) & MULTS_1_2_1(0,3)(PERCISION downto 1));
			MULTS_2_3_1(0,3)<=signed(MULTS_1_3_1(0,3)(PERCISION) & MULTS_1_3_1(0,3)(PERCISION downto 1));
			MULTS_2_4_1(0,3)<=signed(MULTS_1_4_1(0,3)(PERCISION) & MULTS_1_4_1(0,3)(PERCISION downto 1));
			MULTS_2_5_1(0,3)<=signed(MULTS_1_5_1(0,3)(PERCISION) & MULTS_1_5_1(0,3)(PERCISION downto 1));
			MULTS_2_6_1(0,3)<=signed(MULTS_1_6_1(0,3)(PERCISION) & MULTS_1_6_1(0,3)(PERCISION downto 1));
			MULTS_2_7_1(0,3)<=signed(MULTS_1_7_1(0,3)(PERCISION) & MULTS_1_7_1(0,3)(PERCISION downto 1));
			MULTS_2_8_1(0,3)<=signed(MULTS_1_8_1(0,3)(PERCISION) & MULTS_1_8_1(0,3)(PERCISION downto 1));
			MULTS_2_9_1(0,3)<=signed(MULTS_1_9_1(0,3)(PERCISION) & MULTS_1_9_1(0,3)(PERCISION downto 1));
			MULTS_2_10_1(0,3)<=signed(MULTS_1_10_1(0,3)(PERCISION) & MULTS_1_10_1(0,3)(PERCISION downto 1));
			MULTS_2_11_1(0,3)<=signed(MULTS_1_11_1(0,3)(PERCISION) & MULTS_1_11_1(0,3)(PERCISION downto 1));
			MULTS_2_12_1(0,3)<=signed(MULTS_1_12_1(0,3)(PERCISION) & MULTS_1_12_1(0,3)(PERCISION downto 1));
			MULTS_2_13_1(0,3)<=signed(MULTS_1_13_1(0,3)(PERCISION) & MULTS_1_13_1(0,3)(PERCISION downto 1));
			MULTS_2_14_1(0,3)<=signed(MULTS_1_14_1(0,3)(PERCISION) & MULTS_1_14_1(0,3)(PERCISION downto 1));
			MULTS_2_15_1(0,3)<=signed(MULTS_1_15_1(0,3)(PERCISION) & MULTS_1_15_1(0,3)(PERCISION downto 1));
			MULTS_2_16_1(0,3)<=signed(MULTS_1_16_1(0,3)(PERCISION) & MULTS_1_16_1(0,3)(PERCISION downto 1));

			MULTS_2_1_1(0,4)<=signed(MULTS_1_1_1(0,4)(PERCISION) & MULTS_1_1_1(0,4)(PERCISION downto 1));
			MULTS_2_2_1(0,4)<=signed(MULTS_1_2_1(0,4)(PERCISION) & MULTS_1_2_1(0,4)(PERCISION downto 1));
			MULTS_2_3_1(0,4)<=signed(MULTS_1_3_1(0,4)(PERCISION) & MULTS_1_3_1(0,4)(PERCISION downto 1));
			MULTS_2_4_1(0,4)<=signed(MULTS_1_4_1(0,4)(PERCISION) & MULTS_1_4_1(0,4)(PERCISION downto 1));
			MULTS_2_5_1(0,4)<=signed(MULTS_1_5_1(0,4)(PERCISION) & MULTS_1_5_1(0,4)(PERCISION downto 1));
			MULTS_2_6_1(0,4)<=signed(MULTS_1_6_1(0,4)(PERCISION) & MULTS_1_6_1(0,4)(PERCISION downto 1));
			MULTS_2_7_1(0,4)<=signed(MULTS_1_7_1(0,4)(PERCISION) & MULTS_1_7_1(0,4)(PERCISION downto 1));
			MULTS_2_8_1(0,4)<=signed(MULTS_1_8_1(0,4)(PERCISION) & MULTS_1_8_1(0,4)(PERCISION downto 1));
			MULTS_2_9_1(0,4)<=signed(MULTS_1_9_1(0,4)(PERCISION) & MULTS_1_9_1(0,4)(PERCISION downto 1));
			MULTS_2_10_1(0,4)<=signed(MULTS_1_10_1(0,4)(PERCISION) & MULTS_1_10_1(0,4)(PERCISION downto 1));
			MULTS_2_11_1(0,4)<=signed(MULTS_1_11_1(0,4)(PERCISION) & MULTS_1_11_1(0,4)(PERCISION downto 1));
			MULTS_2_12_1(0,4)<=signed(MULTS_1_12_1(0,4)(PERCISION) & MULTS_1_12_1(0,4)(PERCISION downto 1));
			MULTS_2_13_1(0,4)<=signed(MULTS_1_13_1(0,4)(PERCISION) & MULTS_1_13_1(0,4)(PERCISION downto 1));
			MULTS_2_14_1(0,4)<=signed(MULTS_1_14_1(0,4)(PERCISION) & MULTS_1_14_1(0,4)(PERCISION downto 1));
			MULTS_2_15_1(0,4)<=signed(MULTS_1_15_1(0,4)(PERCISION) & MULTS_1_15_1(0,4)(PERCISION downto 1));
			MULTS_2_16_1(0,4)<=signed(MULTS_1_16_1(0,4)(PERCISION) & MULTS_1_16_1(0,4)(PERCISION downto 1));

			MULTS_2_1_1(1,0)<=signed(MULTS_1_1_1(1,0)(PERCISION) & MULTS_1_1_1(1,0)(PERCISION downto 1));
			MULTS_2_2_1(1,0)<=signed(MULTS_1_2_1(1,0)(PERCISION) & MULTS_1_2_1(1,0)(PERCISION downto 1));
			MULTS_2_3_1(1,0)<=signed(MULTS_1_3_1(1,0)(PERCISION) & MULTS_1_3_1(1,0)(PERCISION downto 1));
			MULTS_2_4_1(1,0)<=signed(MULTS_1_4_1(1,0)(PERCISION) & MULTS_1_4_1(1,0)(PERCISION downto 1));
			MULTS_2_5_1(1,0)<=signed(MULTS_1_5_1(1,0)(PERCISION) & MULTS_1_5_1(1,0)(PERCISION downto 1));
			MULTS_2_6_1(1,0)<=signed(MULTS_1_6_1(1,0)(PERCISION) & MULTS_1_6_1(1,0)(PERCISION downto 1));
			MULTS_2_7_1(1,0)<=signed(MULTS_1_7_1(1,0)(PERCISION) & MULTS_1_7_1(1,0)(PERCISION downto 1));
			MULTS_2_8_1(1,0)<=signed(MULTS_1_8_1(1,0)(PERCISION) & MULTS_1_8_1(1,0)(PERCISION downto 1));
			MULTS_2_9_1(1,0)<=signed(MULTS_1_9_1(1,0)(PERCISION) & MULTS_1_9_1(1,0)(PERCISION downto 1));
			MULTS_2_10_1(1,0)<=signed(MULTS_1_10_1(1,0)(PERCISION) & MULTS_1_10_1(1,0)(PERCISION downto 1));
			MULTS_2_11_1(1,0)<=signed(MULTS_1_11_1(1,0)(PERCISION) & MULTS_1_11_1(1,0)(PERCISION downto 1));
			MULTS_2_12_1(1,0)<=signed(MULTS_1_12_1(1,0)(PERCISION) & MULTS_1_12_1(1,0)(PERCISION downto 1));
			MULTS_2_13_1(1,0)<=signed(MULTS_1_13_1(1,0)(PERCISION) & MULTS_1_13_1(1,0)(PERCISION downto 1));
			MULTS_2_14_1(1,0)<=signed(MULTS_1_14_1(1,0)(PERCISION) & MULTS_1_14_1(1,0)(PERCISION downto 1));
			MULTS_2_15_1(1,0)<=signed(MULTS_1_15_1(1,0)(PERCISION) & MULTS_1_15_1(1,0)(PERCISION downto 1));
			MULTS_2_16_1(1,0)<=signed(MULTS_1_16_1(1,0)(PERCISION) & MULTS_1_16_1(1,0)(PERCISION downto 1));

			MULTS_2_1_1(1,1)<=signed(MULTS_1_1_1(1,1)(PERCISION) & MULTS_1_1_1(1,1)(PERCISION downto 1));
			MULTS_2_2_1(1,1)<=signed(MULTS_1_2_1(1,1)(PERCISION) & MULTS_1_2_1(1,1)(PERCISION downto 1));
			MULTS_2_3_1(1,1)<=signed(MULTS_1_3_1(1,1)(PERCISION) & MULTS_1_3_1(1,1)(PERCISION downto 1));
			MULTS_2_4_1(1,1)<=signed(MULTS_1_4_1(1,1)(PERCISION) & MULTS_1_4_1(1,1)(PERCISION downto 1));
			MULTS_2_5_1(1,1)<=signed(MULTS_1_5_1(1,1)(PERCISION) & MULTS_1_5_1(1,1)(PERCISION downto 1));
			MULTS_2_6_1(1,1)<=signed(MULTS_1_6_1(1,1)(PERCISION) & MULTS_1_6_1(1,1)(PERCISION downto 1));
			MULTS_2_7_1(1,1)<=signed(MULTS_1_7_1(1,1)(PERCISION) & MULTS_1_7_1(1,1)(PERCISION downto 1));
			MULTS_2_8_1(1,1)<=signed(MULTS_1_8_1(1,1)(PERCISION) & MULTS_1_8_1(1,1)(PERCISION downto 1));
			MULTS_2_9_1(1,1)<=signed(MULTS_1_9_1(1,1)(PERCISION) & MULTS_1_9_1(1,1)(PERCISION downto 1));
			MULTS_2_10_1(1,1)<=signed(MULTS_1_10_1(1,1)(PERCISION) & MULTS_1_10_1(1,1)(PERCISION downto 1));
			MULTS_2_11_1(1,1)<=signed(MULTS_1_11_1(1,1)(PERCISION) & MULTS_1_11_1(1,1)(PERCISION downto 1));
			MULTS_2_12_1(1,1)<=signed(MULTS_1_12_1(1,1)(PERCISION) & MULTS_1_12_1(1,1)(PERCISION downto 1));
			MULTS_2_13_1(1,1)<=signed(MULTS_1_13_1(1,1)(PERCISION) & MULTS_1_13_1(1,1)(PERCISION downto 1));
			MULTS_2_14_1(1,1)<=signed(MULTS_1_14_1(1,1)(PERCISION) & MULTS_1_14_1(1,1)(PERCISION downto 1));
			MULTS_2_15_1(1,1)<=signed(MULTS_1_15_1(1,1)(PERCISION) & MULTS_1_15_1(1,1)(PERCISION downto 1));
			MULTS_2_16_1(1,1)<=signed(MULTS_1_16_1(1,1)(PERCISION) & MULTS_1_16_1(1,1)(PERCISION downto 1));

			MULTS_2_1_1(1,2)<=signed(MULTS_1_1_1(1,2)(PERCISION) & MULTS_1_1_1(1,2)(PERCISION downto 1));
			MULTS_2_2_1(1,2)<=signed(MULTS_1_2_1(1,2)(PERCISION) & MULTS_1_2_1(1,2)(PERCISION downto 1));
			MULTS_2_3_1(1,2)<=signed(MULTS_1_3_1(1,2)(PERCISION) & MULTS_1_3_1(1,2)(PERCISION downto 1));
			MULTS_2_4_1(1,2)<=signed(MULTS_1_4_1(1,2)(PERCISION) & MULTS_1_4_1(1,2)(PERCISION downto 1));
			MULTS_2_5_1(1,2)<=signed(MULTS_1_5_1(1,2)(PERCISION) & MULTS_1_5_1(1,2)(PERCISION downto 1));
			MULTS_2_6_1(1,2)<=signed(MULTS_1_6_1(1,2)(PERCISION) & MULTS_1_6_1(1,2)(PERCISION downto 1));
			MULTS_2_7_1(1,2)<=signed(MULTS_1_7_1(1,2)(PERCISION) & MULTS_1_7_1(1,2)(PERCISION downto 1));
			MULTS_2_8_1(1,2)<=signed(MULTS_1_8_1(1,2)(PERCISION) & MULTS_1_8_1(1,2)(PERCISION downto 1));
			MULTS_2_9_1(1,2)<=signed(MULTS_1_9_1(1,2)(PERCISION) & MULTS_1_9_1(1,2)(PERCISION downto 1));
			MULTS_2_10_1(1,2)<=signed(MULTS_1_10_1(1,2)(PERCISION) & MULTS_1_10_1(1,2)(PERCISION downto 1));
			MULTS_2_11_1(1,2)<=signed(MULTS_1_11_1(1,2)(PERCISION) & MULTS_1_11_1(1,2)(PERCISION downto 1));
			MULTS_2_12_1(1,2)<=signed(MULTS_1_12_1(1,2)(PERCISION) & MULTS_1_12_1(1,2)(PERCISION downto 1));
			MULTS_2_13_1(1,2)<=signed(MULTS_1_13_1(1,2)(PERCISION) & MULTS_1_13_1(1,2)(PERCISION downto 1));
			MULTS_2_14_1(1,2)<=signed(MULTS_1_14_1(1,2)(PERCISION) & MULTS_1_14_1(1,2)(PERCISION downto 1));
			MULTS_2_15_1(1,2)<=signed(MULTS_1_15_1(1,2)(PERCISION) & MULTS_1_15_1(1,2)(PERCISION downto 1));
			MULTS_2_16_1(1,2)<=signed(MULTS_1_16_1(1,2)(PERCISION) & MULTS_1_16_1(1,2)(PERCISION downto 1));

			MULTS_2_1_1(1,3)<=signed(MULTS_1_1_1(1,3)(PERCISION) & MULTS_1_1_1(1,3)(PERCISION downto 1));
			MULTS_2_2_1(1,3)<=signed(MULTS_1_2_1(1,3)(PERCISION) & MULTS_1_2_1(1,3)(PERCISION downto 1));
			MULTS_2_3_1(1,3)<=signed(MULTS_1_3_1(1,3)(PERCISION) & MULTS_1_3_1(1,3)(PERCISION downto 1));
			MULTS_2_4_1(1,3)<=signed(MULTS_1_4_1(1,3)(PERCISION) & MULTS_1_4_1(1,3)(PERCISION downto 1));
			MULTS_2_5_1(1,3)<=signed(MULTS_1_5_1(1,3)(PERCISION) & MULTS_1_5_1(1,3)(PERCISION downto 1));
			MULTS_2_6_1(1,3)<=signed(MULTS_1_6_1(1,3)(PERCISION) & MULTS_1_6_1(1,3)(PERCISION downto 1));
			MULTS_2_7_1(1,3)<=signed(MULTS_1_7_1(1,3)(PERCISION) & MULTS_1_7_1(1,3)(PERCISION downto 1));
			MULTS_2_8_1(1,3)<=signed(MULTS_1_8_1(1,3)(PERCISION) & MULTS_1_8_1(1,3)(PERCISION downto 1));
			MULTS_2_9_1(1,3)<=signed(MULTS_1_9_1(1,3)(PERCISION) & MULTS_1_9_1(1,3)(PERCISION downto 1));
			MULTS_2_10_1(1,3)<=signed(MULTS_1_10_1(1,3)(PERCISION) & MULTS_1_10_1(1,3)(PERCISION downto 1));
			MULTS_2_11_1(1,3)<=signed(MULTS_1_11_1(1,3)(PERCISION) & MULTS_1_11_1(1,3)(PERCISION downto 1));
			MULTS_2_12_1(1,3)<=signed(MULTS_1_12_1(1,3)(PERCISION) & MULTS_1_12_1(1,3)(PERCISION downto 1));
			MULTS_2_13_1(1,3)<=signed(MULTS_1_13_1(1,3)(PERCISION) & MULTS_1_13_1(1,3)(PERCISION downto 1));
			MULTS_2_14_1(1,3)<=signed(MULTS_1_14_1(1,3)(PERCISION) & MULTS_1_14_1(1,3)(PERCISION downto 1));
			MULTS_2_15_1(1,3)<=signed(MULTS_1_15_1(1,3)(PERCISION) & MULTS_1_15_1(1,3)(PERCISION downto 1));
			MULTS_2_16_1(1,3)<=signed(MULTS_1_16_1(1,3)(PERCISION) & MULTS_1_16_1(1,3)(PERCISION downto 1));

			MULTS_2_1_1(1,4)<=signed(MULTS_1_1_1(1,4)(PERCISION) & MULTS_1_1_1(1,4)(PERCISION downto 1));
			MULTS_2_2_1(1,4)<=signed(MULTS_1_2_1(1,4)(PERCISION) & MULTS_1_2_1(1,4)(PERCISION downto 1));
			MULTS_2_3_1(1,4)<=signed(MULTS_1_3_1(1,4)(PERCISION) & MULTS_1_3_1(1,4)(PERCISION downto 1));
			MULTS_2_4_1(1,4)<=signed(MULTS_1_4_1(1,4)(PERCISION) & MULTS_1_4_1(1,4)(PERCISION downto 1));
			MULTS_2_5_1(1,4)<=signed(MULTS_1_5_1(1,4)(PERCISION) & MULTS_1_5_1(1,4)(PERCISION downto 1));
			MULTS_2_6_1(1,4)<=signed(MULTS_1_6_1(1,4)(PERCISION) & MULTS_1_6_1(1,4)(PERCISION downto 1));
			MULTS_2_7_1(1,4)<=signed(MULTS_1_7_1(1,4)(PERCISION) & MULTS_1_7_1(1,4)(PERCISION downto 1));
			MULTS_2_8_1(1,4)<=signed(MULTS_1_8_1(1,4)(PERCISION) & MULTS_1_8_1(1,4)(PERCISION downto 1));
			MULTS_2_9_1(1,4)<=signed(MULTS_1_9_1(1,4)(PERCISION) & MULTS_1_9_1(1,4)(PERCISION downto 1));
			MULTS_2_10_1(1,4)<=signed(MULTS_1_10_1(1,4)(PERCISION) & MULTS_1_10_1(1,4)(PERCISION downto 1));
			MULTS_2_11_1(1,4)<=signed(MULTS_1_11_1(1,4)(PERCISION) & MULTS_1_11_1(1,4)(PERCISION downto 1));
			MULTS_2_12_1(1,4)<=signed(MULTS_1_12_1(1,4)(PERCISION) & MULTS_1_12_1(1,4)(PERCISION downto 1));
			MULTS_2_13_1(1,4)<=signed(MULTS_1_13_1(1,4)(PERCISION) & MULTS_1_13_1(1,4)(PERCISION downto 1));
			MULTS_2_14_1(1,4)<=signed(MULTS_1_14_1(1,4)(PERCISION) & MULTS_1_14_1(1,4)(PERCISION downto 1));
			MULTS_2_15_1(1,4)<=signed(MULTS_1_15_1(1,4)(PERCISION) & MULTS_1_15_1(1,4)(PERCISION downto 1));
			MULTS_2_16_1(1,4)<=signed(MULTS_1_16_1(1,4)(PERCISION) & MULTS_1_16_1(1,4)(PERCISION downto 1));

			MULTS_2_1_1(2,0)<=signed(MULTS_1_1_1(2,0)(PERCISION) & MULTS_1_1_1(2,0)(PERCISION downto 1));
			MULTS_2_2_1(2,0)<=signed(MULTS_1_2_1(2,0)(PERCISION) & MULTS_1_2_1(2,0)(PERCISION downto 1));
			MULTS_2_3_1(2,0)<=signed(MULTS_1_3_1(2,0)(PERCISION) & MULTS_1_3_1(2,0)(PERCISION downto 1));
			MULTS_2_4_1(2,0)<=signed(MULTS_1_4_1(2,0)(PERCISION) & MULTS_1_4_1(2,0)(PERCISION downto 1));
			MULTS_2_5_1(2,0)<=signed(MULTS_1_5_1(2,0)(PERCISION) & MULTS_1_5_1(2,0)(PERCISION downto 1));
			MULTS_2_6_1(2,0)<=signed(MULTS_1_6_1(2,0)(PERCISION) & MULTS_1_6_1(2,0)(PERCISION downto 1));
			MULTS_2_7_1(2,0)<=signed(MULTS_1_7_1(2,0)(PERCISION) & MULTS_1_7_1(2,0)(PERCISION downto 1));
			MULTS_2_8_1(2,0)<=signed(MULTS_1_8_1(2,0)(PERCISION) & MULTS_1_8_1(2,0)(PERCISION downto 1));
			MULTS_2_9_1(2,0)<=signed(MULTS_1_9_1(2,0)(PERCISION) & MULTS_1_9_1(2,0)(PERCISION downto 1));
			MULTS_2_10_1(2,0)<=signed(MULTS_1_10_1(2,0)(PERCISION) & MULTS_1_10_1(2,0)(PERCISION downto 1));
			MULTS_2_11_1(2,0)<=signed(MULTS_1_11_1(2,0)(PERCISION) & MULTS_1_11_1(2,0)(PERCISION downto 1));
			MULTS_2_12_1(2,0)<=signed(MULTS_1_12_1(2,0)(PERCISION) & MULTS_1_12_1(2,0)(PERCISION downto 1));
			MULTS_2_13_1(2,0)<=signed(MULTS_1_13_1(2,0)(PERCISION) & MULTS_1_13_1(2,0)(PERCISION downto 1));
			MULTS_2_14_1(2,0)<=signed(MULTS_1_14_1(2,0)(PERCISION) & MULTS_1_14_1(2,0)(PERCISION downto 1));
			MULTS_2_15_1(2,0)<=signed(MULTS_1_15_1(2,0)(PERCISION) & MULTS_1_15_1(2,0)(PERCISION downto 1));
			MULTS_2_16_1(2,0)<=signed(MULTS_1_16_1(2,0)(PERCISION) & MULTS_1_16_1(2,0)(PERCISION downto 1));

			MULTS_2_1_1(2,1)<=signed(MULTS_1_1_1(2,1)(PERCISION) & MULTS_1_1_1(2,1)(PERCISION downto 1));
			MULTS_2_2_1(2,1)<=signed(MULTS_1_2_1(2,1)(PERCISION) & MULTS_1_2_1(2,1)(PERCISION downto 1));
			MULTS_2_3_1(2,1)<=signed(MULTS_1_3_1(2,1)(PERCISION) & MULTS_1_3_1(2,1)(PERCISION downto 1));
			MULTS_2_4_1(2,1)<=signed(MULTS_1_4_1(2,1)(PERCISION) & MULTS_1_4_1(2,1)(PERCISION downto 1));
			MULTS_2_5_1(2,1)<=signed(MULTS_1_5_1(2,1)(PERCISION) & MULTS_1_5_1(2,1)(PERCISION downto 1));
			MULTS_2_6_1(2,1)<=signed(MULTS_1_6_1(2,1)(PERCISION) & MULTS_1_6_1(2,1)(PERCISION downto 1));
			MULTS_2_7_1(2,1)<=signed(MULTS_1_7_1(2,1)(PERCISION) & MULTS_1_7_1(2,1)(PERCISION downto 1));
			MULTS_2_8_1(2,1)<=signed(MULTS_1_8_1(2,1)(PERCISION) & MULTS_1_8_1(2,1)(PERCISION downto 1));
			MULTS_2_9_1(2,1)<=signed(MULTS_1_9_1(2,1)(PERCISION) & MULTS_1_9_1(2,1)(PERCISION downto 1));
			MULTS_2_10_1(2,1)<=signed(MULTS_1_10_1(2,1)(PERCISION) & MULTS_1_10_1(2,1)(PERCISION downto 1));
			MULTS_2_11_1(2,1)<=signed(MULTS_1_11_1(2,1)(PERCISION) & MULTS_1_11_1(2,1)(PERCISION downto 1));
			MULTS_2_12_1(2,1)<=signed(MULTS_1_12_1(2,1)(PERCISION) & MULTS_1_12_1(2,1)(PERCISION downto 1));
			MULTS_2_13_1(2,1)<=signed(MULTS_1_13_1(2,1)(PERCISION) & MULTS_1_13_1(2,1)(PERCISION downto 1));
			MULTS_2_14_1(2,1)<=signed(MULTS_1_14_1(2,1)(PERCISION) & MULTS_1_14_1(2,1)(PERCISION downto 1));
			MULTS_2_15_1(2,1)<=signed(MULTS_1_15_1(2,1)(PERCISION) & MULTS_1_15_1(2,1)(PERCISION downto 1));
			MULTS_2_16_1(2,1)<=signed(MULTS_1_16_1(2,1)(PERCISION) & MULTS_1_16_1(2,1)(PERCISION downto 1));

			MULTS_2_1_1(2,2)<=signed(MULTS_1_1_1(2,2)(PERCISION) & MULTS_1_1_1(2,2)(PERCISION downto 1));
			MULTS_2_2_1(2,2)<=signed(MULTS_1_2_1(2,2)(PERCISION) & MULTS_1_2_1(2,2)(PERCISION downto 1));
			MULTS_2_3_1(2,2)<=signed(MULTS_1_3_1(2,2)(PERCISION) & MULTS_1_3_1(2,2)(PERCISION downto 1));
			MULTS_2_4_1(2,2)<=signed(MULTS_1_4_1(2,2)(PERCISION) & MULTS_1_4_1(2,2)(PERCISION downto 1));
			MULTS_2_5_1(2,2)<=signed(MULTS_1_5_1(2,2)(PERCISION) & MULTS_1_5_1(2,2)(PERCISION downto 1));
			MULTS_2_6_1(2,2)<=signed(MULTS_1_6_1(2,2)(PERCISION) & MULTS_1_6_1(2,2)(PERCISION downto 1));
			MULTS_2_7_1(2,2)<=signed(MULTS_1_7_1(2,2)(PERCISION) & MULTS_1_7_1(2,2)(PERCISION downto 1));
			MULTS_2_8_1(2,2)<=signed(MULTS_1_8_1(2,2)(PERCISION) & MULTS_1_8_1(2,2)(PERCISION downto 1));
			MULTS_2_9_1(2,2)<=signed(MULTS_1_9_1(2,2)(PERCISION) & MULTS_1_9_1(2,2)(PERCISION downto 1));
			MULTS_2_10_1(2,2)<=signed(MULTS_1_10_1(2,2)(PERCISION) & MULTS_1_10_1(2,2)(PERCISION downto 1));
			MULTS_2_11_1(2,2)<=signed(MULTS_1_11_1(2,2)(PERCISION) & MULTS_1_11_1(2,2)(PERCISION downto 1));
			MULTS_2_12_1(2,2)<=signed(MULTS_1_12_1(2,2)(PERCISION) & MULTS_1_12_1(2,2)(PERCISION downto 1));
			MULTS_2_13_1(2,2)<=signed(MULTS_1_13_1(2,2)(PERCISION) & MULTS_1_13_1(2,2)(PERCISION downto 1));
			MULTS_2_14_1(2,2)<=signed(MULTS_1_14_1(2,2)(PERCISION) & MULTS_1_14_1(2,2)(PERCISION downto 1));
			MULTS_2_15_1(2,2)<=signed(MULTS_1_15_1(2,2)(PERCISION) & MULTS_1_15_1(2,2)(PERCISION downto 1));
			MULTS_2_16_1(2,2)<=signed(MULTS_1_16_1(2,2)(PERCISION) & MULTS_1_16_1(2,2)(PERCISION downto 1));

			MULTS_2_1_1(2,3)<=signed(MULTS_1_1_1(2,3)(PERCISION) & MULTS_1_1_1(2,3)(PERCISION downto 1));
			MULTS_2_2_1(2,3)<=signed(MULTS_1_2_1(2,3)(PERCISION) & MULTS_1_2_1(2,3)(PERCISION downto 1));
			MULTS_2_3_1(2,3)<=signed(MULTS_1_3_1(2,3)(PERCISION) & MULTS_1_3_1(2,3)(PERCISION downto 1));
			MULTS_2_4_1(2,3)<=signed(MULTS_1_4_1(2,3)(PERCISION) & MULTS_1_4_1(2,3)(PERCISION downto 1));
			MULTS_2_5_1(2,3)<=signed(MULTS_1_5_1(2,3)(PERCISION) & MULTS_1_5_1(2,3)(PERCISION downto 1));
			MULTS_2_6_1(2,3)<=signed(MULTS_1_6_1(2,3)(PERCISION) & MULTS_1_6_1(2,3)(PERCISION downto 1));
			MULTS_2_7_1(2,3)<=signed(MULTS_1_7_1(2,3)(PERCISION) & MULTS_1_7_1(2,3)(PERCISION downto 1));
			MULTS_2_8_1(2,3)<=signed(MULTS_1_8_1(2,3)(PERCISION) & MULTS_1_8_1(2,3)(PERCISION downto 1));
			MULTS_2_9_1(2,3)<=signed(MULTS_1_9_1(2,3)(PERCISION) & MULTS_1_9_1(2,3)(PERCISION downto 1));
			MULTS_2_10_1(2,3)<=signed(MULTS_1_10_1(2,3)(PERCISION) & MULTS_1_10_1(2,3)(PERCISION downto 1));
			MULTS_2_11_1(2,3)<=signed(MULTS_1_11_1(2,3)(PERCISION) & MULTS_1_11_1(2,3)(PERCISION downto 1));
			MULTS_2_12_1(2,3)<=signed(MULTS_1_12_1(2,3)(PERCISION) & MULTS_1_12_1(2,3)(PERCISION downto 1));
			MULTS_2_13_1(2,3)<=signed(MULTS_1_13_1(2,3)(PERCISION) & MULTS_1_13_1(2,3)(PERCISION downto 1));
			MULTS_2_14_1(2,3)<=signed(MULTS_1_14_1(2,3)(PERCISION) & MULTS_1_14_1(2,3)(PERCISION downto 1));
			MULTS_2_15_1(2,3)<=signed(MULTS_1_15_1(2,3)(PERCISION) & MULTS_1_15_1(2,3)(PERCISION downto 1));
			MULTS_2_16_1(2,3)<=signed(MULTS_1_16_1(2,3)(PERCISION) & MULTS_1_16_1(2,3)(PERCISION downto 1));

			MULTS_2_1_1(2,4)<=signed(MULTS_1_1_1(2,4)(PERCISION) & MULTS_1_1_1(2,4)(PERCISION downto 1));
			MULTS_2_2_1(2,4)<=signed(MULTS_1_2_1(2,4)(PERCISION) & MULTS_1_2_1(2,4)(PERCISION downto 1));
			MULTS_2_3_1(2,4)<=signed(MULTS_1_3_1(2,4)(PERCISION) & MULTS_1_3_1(2,4)(PERCISION downto 1));
			MULTS_2_4_1(2,4)<=signed(MULTS_1_4_1(2,4)(PERCISION) & MULTS_1_4_1(2,4)(PERCISION downto 1));
			MULTS_2_5_1(2,4)<=signed(MULTS_1_5_1(2,4)(PERCISION) & MULTS_1_5_1(2,4)(PERCISION downto 1));
			MULTS_2_6_1(2,4)<=signed(MULTS_1_6_1(2,4)(PERCISION) & MULTS_1_6_1(2,4)(PERCISION downto 1));
			MULTS_2_7_1(2,4)<=signed(MULTS_1_7_1(2,4)(PERCISION) & MULTS_1_7_1(2,4)(PERCISION downto 1));
			MULTS_2_8_1(2,4)<=signed(MULTS_1_8_1(2,4)(PERCISION) & MULTS_1_8_1(2,4)(PERCISION downto 1));
			MULTS_2_9_1(2,4)<=signed(MULTS_1_9_1(2,4)(PERCISION) & MULTS_1_9_1(2,4)(PERCISION downto 1));
			MULTS_2_10_1(2,4)<=signed(MULTS_1_10_1(2,4)(PERCISION) & MULTS_1_10_1(2,4)(PERCISION downto 1));
			MULTS_2_11_1(2,4)<=signed(MULTS_1_11_1(2,4)(PERCISION) & MULTS_1_11_1(2,4)(PERCISION downto 1));
			MULTS_2_12_1(2,4)<=signed(MULTS_1_12_1(2,4)(PERCISION) & MULTS_1_12_1(2,4)(PERCISION downto 1));
			MULTS_2_13_1(2,4)<=signed(MULTS_1_13_1(2,4)(PERCISION) & MULTS_1_13_1(2,4)(PERCISION downto 1));
			MULTS_2_14_1(2,4)<=signed(MULTS_1_14_1(2,4)(PERCISION) & MULTS_1_14_1(2,4)(PERCISION downto 1));
			MULTS_2_15_1(2,4)<=signed(MULTS_1_15_1(2,4)(PERCISION) & MULTS_1_15_1(2,4)(PERCISION downto 1));
			MULTS_2_16_1(2,4)<=signed(MULTS_1_16_1(2,4)(PERCISION) & MULTS_1_16_1(2,4)(PERCISION downto 1));

			MULTS_2_1_1(3,0)<=signed(MULTS_1_1_1(3,0)(PERCISION) & MULTS_1_1_1(3,0)(PERCISION downto 1));
			MULTS_2_2_1(3,0)<=signed(MULTS_1_2_1(3,0)(PERCISION) & MULTS_1_2_1(3,0)(PERCISION downto 1));
			MULTS_2_3_1(3,0)<=signed(MULTS_1_3_1(3,0)(PERCISION) & MULTS_1_3_1(3,0)(PERCISION downto 1));
			MULTS_2_4_1(3,0)<=signed(MULTS_1_4_1(3,0)(PERCISION) & MULTS_1_4_1(3,0)(PERCISION downto 1));
			MULTS_2_5_1(3,0)<=signed(MULTS_1_5_1(3,0)(PERCISION) & MULTS_1_5_1(3,0)(PERCISION downto 1));
			MULTS_2_6_1(3,0)<=signed(MULTS_1_6_1(3,0)(PERCISION) & MULTS_1_6_1(3,0)(PERCISION downto 1));
			MULTS_2_7_1(3,0)<=signed(MULTS_1_7_1(3,0)(PERCISION) & MULTS_1_7_1(3,0)(PERCISION downto 1));
			MULTS_2_8_1(3,0)<=signed(MULTS_1_8_1(3,0)(PERCISION) & MULTS_1_8_1(3,0)(PERCISION downto 1));
			MULTS_2_9_1(3,0)<=signed(MULTS_1_9_1(3,0)(PERCISION) & MULTS_1_9_1(3,0)(PERCISION downto 1));
			MULTS_2_10_1(3,0)<=signed(MULTS_1_10_1(3,0)(PERCISION) & MULTS_1_10_1(3,0)(PERCISION downto 1));
			MULTS_2_11_1(3,0)<=signed(MULTS_1_11_1(3,0)(PERCISION) & MULTS_1_11_1(3,0)(PERCISION downto 1));
			MULTS_2_12_1(3,0)<=signed(MULTS_1_12_1(3,0)(PERCISION) & MULTS_1_12_1(3,0)(PERCISION downto 1));
			MULTS_2_13_1(3,0)<=signed(MULTS_1_13_1(3,0)(PERCISION) & MULTS_1_13_1(3,0)(PERCISION downto 1));
			MULTS_2_14_1(3,0)<=signed(MULTS_1_14_1(3,0)(PERCISION) & MULTS_1_14_1(3,0)(PERCISION downto 1));
			MULTS_2_15_1(3,0)<=signed(MULTS_1_15_1(3,0)(PERCISION) & MULTS_1_15_1(3,0)(PERCISION downto 1));
			MULTS_2_16_1(3,0)<=signed(MULTS_1_16_1(3,0)(PERCISION) & MULTS_1_16_1(3,0)(PERCISION downto 1));

			MULTS_2_1_1(3,1)<=signed(MULTS_1_1_1(3,1)(PERCISION) & MULTS_1_1_1(3,1)(PERCISION downto 1));
			MULTS_2_2_1(3,1)<=signed(MULTS_1_2_1(3,1)(PERCISION) & MULTS_1_2_1(3,1)(PERCISION downto 1));
			MULTS_2_3_1(3,1)<=signed(MULTS_1_3_1(3,1)(PERCISION) & MULTS_1_3_1(3,1)(PERCISION downto 1));
			MULTS_2_4_1(3,1)<=signed(MULTS_1_4_1(3,1)(PERCISION) & MULTS_1_4_1(3,1)(PERCISION downto 1));
			MULTS_2_5_1(3,1)<=signed(MULTS_1_5_1(3,1)(PERCISION) & MULTS_1_5_1(3,1)(PERCISION downto 1));
			MULTS_2_6_1(3,1)<=signed(MULTS_1_6_1(3,1)(PERCISION) & MULTS_1_6_1(3,1)(PERCISION downto 1));
			MULTS_2_7_1(3,1)<=signed(MULTS_1_7_1(3,1)(PERCISION) & MULTS_1_7_1(3,1)(PERCISION downto 1));
			MULTS_2_8_1(3,1)<=signed(MULTS_1_8_1(3,1)(PERCISION) & MULTS_1_8_1(3,1)(PERCISION downto 1));
			MULTS_2_9_1(3,1)<=signed(MULTS_1_9_1(3,1)(PERCISION) & MULTS_1_9_1(3,1)(PERCISION downto 1));
			MULTS_2_10_1(3,1)<=signed(MULTS_1_10_1(3,1)(PERCISION) & MULTS_1_10_1(3,1)(PERCISION downto 1));
			MULTS_2_11_1(3,1)<=signed(MULTS_1_11_1(3,1)(PERCISION) & MULTS_1_11_1(3,1)(PERCISION downto 1));
			MULTS_2_12_1(3,1)<=signed(MULTS_1_12_1(3,1)(PERCISION) & MULTS_1_12_1(3,1)(PERCISION downto 1));
			MULTS_2_13_1(3,1)<=signed(MULTS_1_13_1(3,1)(PERCISION) & MULTS_1_13_1(3,1)(PERCISION downto 1));
			MULTS_2_14_1(3,1)<=signed(MULTS_1_14_1(3,1)(PERCISION) & MULTS_1_14_1(3,1)(PERCISION downto 1));
			MULTS_2_15_1(3,1)<=signed(MULTS_1_15_1(3,1)(PERCISION) & MULTS_1_15_1(3,1)(PERCISION downto 1));
			MULTS_2_16_1(3,1)<=signed(MULTS_1_16_1(3,1)(PERCISION) & MULTS_1_16_1(3,1)(PERCISION downto 1));

			MULTS_2_1_1(3,2)<=signed(MULTS_1_1_1(3,2)(PERCISION) & MULTS_1_1_1(3,2)(PERCISION downto 1));
			MULTS_2_2_1(3,2)<=signed(MULTS_1_2_1(3,2)(PERCISION) & MULTS_1_2_1(3,2)(PERCISION downto 1));
			MULTS_2_3_1(3,2)<=signed(MULTS_1_3_1(3,2)(PERCISION) & MULTS_1_3_1(3,2)(PERCISION downto 1));
			MULTS_2_4_1(3,2)<=signed(MULTS_1_4_1(3,2)(PERCISION) & MULTS_1_4_1(3,2)(PERCISION downto 1));
			MULTS_2_5_1(3,2)<=signed(MULTS_1_5_1(3,2)(PERCISION) & MULTS_1_5_1(3,2)(PERCISION downto 1));
			MULTS_2_6_1(3,2)<=signed(MULTS_1_6_1(3,2)(PERCISION) & MULTS_1_6_1(3,2)(PERCISION downto 1));
			MULTS_2_7_1(3,2)<=signed(MULTS_1_7_1(3,2)(PERCISION) & MULTS_1_7_1(3,2)(PERCISION downto 1));
			MULTS_2_8_1(3,2)<=signed(MULTS_1_8_1(3,2)(PERCISION) & MULTS_1_8_1(3,2)(PERCISION downto 1));
			MULTS_2_9_1(3,2)<=signed(MULTS_1_9_1(3,2)(PERCISION) & MULTS_1_9_1(3,2)(PERCISION downto 1));
			MULTS_2_10_1(3,2)<=signed(MULTS_1_10_1(3,2)(PERCISION) & MULTS_1_10_1(3,2)(PERCISION downto 1));
			MULTS_2_11_1(3,2)<=signed(MULTS_1_11_1(3,2)(PERCISION) & MULTS_1_11_1(3,2)(PERCISION downto 1));
			MULTS_2_12_1(3,2)<=signed(MULTS_1_12_1(3,2)(PERCISION) & MULTS_1_12_1(3,2)(PERCISION downto 1));
			MULTS_2_13_1(3,2)<=signed(MULTS_1_13_1(3,2)(PERCISION) & MULTS_1_13_1(3,2)(PERCISION downto 1));
			MULTS_2_14_1(3,2)<=signed(MULTS_1_14_1(3,2)(PERCISION) & MULTS_1_14_1(3,2)(PERCISION downto 1));
			MULTS_2_15_1(3,2)<=signed(MULTS_1_15_1(3,2)(PERCISION) & MULTS_1_15_1(3,2)(PERCISION downto 1));
			MULTS_2_16_1(3,2)<=signed(MULTS_1_16_1(3,2)(PERCISION) & MULTS_1_16_1(3,2)(PERCISION downto 1));

			MULTS_2_1_1(3,3)<=signed(MULTS_1_1_1(3,3)(PERCISION) & MULTS_1_1_1(3,3)(PERCISION downto 1));
			MULTS_2_2_1(3,3)<=signed(MULTS_1_2_1(3,3)(PERCISION) & MULTS_1_2_1(3,3)(PERCISION downto 1));
			MULTS_2_3_1(3,3)<=signed(MULTS_1_3_1(3,3)(PERCISION) & MULTS_1_3_1(3,3)(PERCISION downto 1));
			MULTS_2_4_1(3,3)<=signed(MULTS_1_4_1(3,3)(PERCISION) & MULTS_1_4_1(3,3)(PERCISION downto 1));
			MULTS_2_5_1(3,3)<=signed(MULTS_1_5_1(3,3)(PERCISION) & MULTS_1_5_1(3,3)(PERCISION downto 1));
			MULTS_2_6_1(3,3)<=signed(MULTS_1_6_1(3,3)(PERCISION) & MULTS_1_6_1(3,3)(PERCISION downto 1));
			MULTS_2_7_1(3,3)<=signed(MULTS_1_7_1(3,3)(PERCISION) & MULTS_1_7_1(3,3)(PERCISION downto 1));
			MULTS_2_8_1(3,3)<=signed(MULTS_1_8_1(3,3)(PERCISION) & MULTS_1_8_1(3,3)(PERCISION downto 1));
			MULTS_2_9_1(3,3)<=signed(MULTS_1_9_1(3,3)(PERCISION) & MULTS_1_9_1(3,3)(PERCISION downto 1));
			MULTS_2_10_1(3,3)<=signed(MULTS_1_10_1(3,3)(PERCISION) & MULTS_1_10_1(3,3)(PERCISION downto 1));
			MULTS_2_11_1(3,3)<=signed(MULTS_1_11_1(3,3)(PERCISION) & MULTS_1_11_1(3,3)(PERCISION downto 1));
			MULTS_2_12_1(3,3)<=signed(MULTS_1_12_1(3,3)(PERCISION) & MULTS_1_12_1(3,3)(PERCISION downto 1));
			MULTS_2_13_1(3,3)<=signed(MULTS_1_13_1(3,3)(PERCISION) & MULTS_1_13_1(3,3)(PERCISION downto 1));
			MULTS_2_14_1(3,3)<=signed(MULTS_1_14_1(3,3)(PERCISION) & MULTS_1_14_1(3,3)(PERCISION downto 1));
			MULTS_2_15_1(3,3)<=signed(MULTS_1_15_1(3,3)(PERCISION) & MULTS_1_15_1(3,3)(PERCISION downto 1));
			MULTS_2_16_1(3,3)<=signed(MULTS_1_16_1(3,3)(PERCISION) & MULTS_1_16_1(3,3)(PERCISION downto 1));

			MULTS_2_1_1(3,4)<=signed(MULTS_1_1_1(3,4)(PERCISION) & MULTS_1_1_1(3,4)(PERCISION downto 1));
			MULTS_2_2_1(3,4)<=signed(MULTS_1_2_1(3,4)(PERCISION) & MULTS_1_2_1(3,4)(PERCISION downto 1));
			MULTS_2_3_1(3,4)<=signed(MULTS_1_3_1(3,4)(PERCISION) & MULTS_1_3_1(3,4)(PERCISION downto 1));
			MULTS_2_4_1(3,4)<=signed(MULTS_1_4_1(3,4)(PERCISION) & MULTS_1_4_1(3,4)(PERCISION downto 1));
			MULTS_2_5_1(3,4)<=signed(MULTS_1_5_1(3,4)(PERCISION) & MULTS_1_5_1(3,4)(PERCISION downto 1));
			MULTS_2_6_1(3,4)<=signed(MULTS_1_6_1(3,4)(PERCISION) & MULTS_1_6_1(3,4)(PERCISION downto 1));
			MULTS_2_7_1(3,4)<=signed(MULTS_1_7_1(3,4)(PERCISION) & MULTS_1_7_1(3,4)(PERCISION downto 1));
			MULTS_2_8_1(3,4)<=signed(MULTS_1_8_1(3,4)(PERCISION) & MULTS_1_8_1(3,4)(PERCISION downto 1));
			MULTS_2_9_1(3,4)<=signed(MULTS_1_9_1(3,4)(PERCISION) & MULTS_1_9_1(3,4)(PERCISION downto 1));
			MULTS_2_10_1(3,4)<=signed(MULTS_1_10_1(3,4)(PERCISION) & MULTS_1_10_1(3,4)(PERCISION downto 1));
			MULTS_2_11_1(3,4)<=signed(MULTS_1_11_1(3,4)(PERCISION) & MULTS_1_11_1(3,4)(PERCISION downto 1));
			MULTS_2_12_1(3,4)<=signed(MULTS_1_12_1(3,4)(PERCISION) & MULTS_1_12_1(3,4)(PERCISION downto 1));
			MULTS_2_13_1(3,4)<=signed(MULTS_1_13_1(3,4)(PERCISION) & MULTS_1_13_1(3,4)(PERCISION downto 1));
			MULTS_2_14_1(3,4)<=signed(MULTS_1_14_1(3,4)(PERCISION) & MULTS_1_14_1(3,4)(PERCISION downto 1));
			MULTS_2_15_1(3,4)<=signed(MULTS_1_15_1(3,4)(PERCISION) & MULTS_1_15_1(3,4)(PERCISION downto 1));
			MULTS_2_16_1(3,4)<=signed(MULTS_1_16_1(3,4)(PERCISION) & MULTS_1_16_1(3,4)(PERCISION downto 1));

			MULTS_2_1_1(4,0)<=signed(MULTS_1_1_1(4,0)(PERCISION) & MULTS_1_1_1(4,0)(PERCISION downto 1));
			MULTS_2_2_1(4,0)<=signed(MULTS_1_2_1(4,0)(PERCISION) & MULTS_1_2_1(4,0)(PERCISION downto 1));
			MULTS_2_3_1(4,0)<=signed(MULTS_1_3_1(4,0)(PERCISION) & MULTS_1_3_1(4,0)(PERCISION downto 1));
			MULTS_2_4_1(4,0)<=signed(MULTS_1_4_1(4,0)(PERCISION) & MULTS_1_4_1(4,0)(PERCISION downto 1));
			MULTS_2_5_1(4,0)<=signed(MULTS_1_5_1(4,0)(PERCISION) & MULTS_1_5_1(4,0)(PERCISION downto 1));
			MULTS_2_6_1(4,0)<=signed(MULTS_1_6_1(4,0)(PERCISION) & MULTS_1_6_1(4,0)(PERCISION downto 1));
			MULTS_2_7_1(4,0)<=signed(MULTS_1_7_1(4,0)(PERCISION) & MULTS_1_7_1(4,0)(PERCISION downto 1));
			MULTS_2_8_1(4,0)<=signed(MULTS_1_8_1(4,0)(PERCISION) & MULTS_1_8_1(4,0)(PERCISION downto 1));
			MULTS_2_9_1(4,0)<=signed(MULTS_1_9_1(4,0)(PERCISION) & MULTS_1_9_1(4,0)(PERCISION downto 1));
			MULTS_2_10_1(4,0)<=signed(MULTS_1_10_1(4,0)(PERCISION) & MULTS_1_10_1(4,0)(PERCISION downto 1));
			MULTS_2_11_1(4,0)<=signed(MULTS_1_11_1(4,0)(PERCISION) & MULTS_1_11_1(4,0)(PERCISION downto 1));
			MULTS_2_12_1(4,0)<=signed(MULTS_1_12_1(4,0)(PERCISION) & MULTS_1_12_1(4,0)(PERCISION downto 1));
			MULTS_2_13_1(4,0)<=signed(MULTS_1_13_1(4,0)(PERCISION) & MULTS_1_13_1(4,0)(PERCISION downto 1));
			MULTS_2_14_1(4,0)<=signed(MULTS_1_14_1(4,0)(PERCISION) & MULTS_1_14_1(4,0)(PERCISION downto 1));
			MULTS_2_15_1(4,0)<=signed(MULTS_1_15_1(4,0)(PERCISION) & MULTS_1_15_1(4,0)(PERCISION downto 1));
			MULTS_2_16_1(4,0)<=signed(MULTS_1_16_1(4,0)(PERCISION) & MULTS_1_16_1(4,0)(PERCISION downto 1));

			MULTS_2_1_1(4,1)<=signed(MULTS_1_1_1(4,1)(PERCISION) & MULTS_1_1_1(4,1)(PERCISION downto 1));
			MULTS_2_2_1(4,1)<=signed(MULTS_1_2_1(4,1)(PERCISION) & MULTS_1_2_1(4,1)(PERCISION downto 1));
			MULTS_2_3_1(4,1)<=signed(MULTS_1_3_1(4,1)(PERCISION) & MULTS_1_3_1(4,1)(PERCISION downto 1));
			MULTS_2_4_1(4,1)<=signed(MULTS_1_4_1(4,1)(PERCISION) & MULTS_1_4_1(4,1)(PERCISION downto 1));
			MULTS_2_5_1(4,1)<=signed(MULTS_1_5_1(4,1)(PERCISION) & MULTS_1_5_1(4,1)(PERCISION downto 1));
			MULTS_2_6_1(4,1)<=signed(MULTS_1_6_1(4,1)(PERCISION) & MULTS_1_6_1(4,1)(PERCISION downto 1));
			MULTS_2_7_1(4,1)<=signed(MULTS_1_7_1(4,1)(PERCISION) & MULTS_1_7_1(4,1)(PERCISION downto 1));
			MULTS_2_8_1(4,1)<=signed(MULTS_1_8_1(4,1)(PERCISION) & MULTS_1_8_1(4,1)(PERCISION downto 1));
			MULTS_2_9_1(4,1)<=signed(MULTS_1_9_1(4,1)(PERCISION) & MULTS_1_9_1(4,1)(PERCISION downto 1));
			MULTS_2_10_1(4,1)<=signed(MULTS_1_10_1(4,1)(PERCISION) & MULTS_1_10_1(4,1)(PERCISION downto 1));
			MULTS_2_11_1(4,1)<=signed(MULTS_1_11_1(4,1)(PERCISION) & MULTS_1_11_1(4,1)(PERCISION downto 1));
			MULTS_2_12_1(4,1)<=signed(MULTS_1_12_1(4,1)(PERCISION) & MULTS_1_12_1(4,1)(PERCISION downto 1));
			MULTS_2_13_1(4,1)<=signed(MULTS_1_13_1(4,1)(PERCISION) & MULTS_1_13_1(4,1)(PERCISION downto 1));
			MULTS_2_14_1(4,1)<=signed(MULTS_1_14_1(4,1)(PERCISION) & MULTS_1_14_1(4,1)(PERCISION downto 1));
			MULTS_2_15_1(4,1)<=signed(MULTS_1_15_1(4,1)(PERCISION) & MULTS_1_15_1(4,1)(PERCISION downto 1));
			MULTS_2_16_1(4,1)<=signed(MULTS_1_16_1(4,1)(PERCISION) & MULTS_1_16_1(4,1)(PERCISION downto 1));

			MULTS_2_1_1(4,2)<=signed(MULTS_1_1_1(4,2)(PERCISION) & MULTS_1_1_1(4,2)(PERCISION downto 1));
			MULTS_2_2_1(4,2)<=signed(MULTS_1_2_1(4,2)(PERCISION) & MULTS_1_2_1(4,2)(PERCISION downto 1));
			MULTS_2_3_1(4,2)<=signed(MULTS_1_3_1(4,2)(PERCISION) & MULTS_1_3_1(4,2)(PERCISION downto 1));
			MULTS_2_4_1(4,2)<=signed(MULTS_1_4_1(4,2)(PERCISION) & MULTS_1_4_1(4,2)(PERCISION downto 1));
			MULTS_2_5_1(4,2)<=signed(MULTS_1_5_1(4,2)(PERCISION) & MULTS_1_5_1(4,2)(PERCISION downto 1));
			MULTS_2_6_1(4,2)<=signed(MULTS_1_6_1(4,2)(PERCISION) & MULTS_1_6_1(4,2)(PERCISION downto 1));
			MULTS_2_7_1(4,2)<=signed(MULTS_1_7_1(4,2)(PERCISION) & MULTS_1_7_1(4,2)(PERCISION downto 1));
			MULTS_2_8_1(4,2)<=signed(MULTS_1_8_1(4,2)(PERCISION) & MULTS_1_8_1(4,2)(PERCISION downto 1));
			MULTS_2_9_1(4,2)<=signed(MULTS_1_9_1(4,2)(PERCISION) & MULTS_1_9_1(4,2)(PERCISION downto 1));
			MULTS_2_10_1(4,2)<=signed(MULTS_1_10_1(4,2)(PERCISION) & MULTS_1_10_1(4,2)(PERCISION downto 1));
			MULTS_2_11_1(4,2)<=signed(MULTS_1_11_1(4,2)(PERCISION) & MULTS_1_11_1(4,2)(PERCISION downto 1));
			MULTS_2_12_1(4,2)<=signed(MULTS_1_12_1(4,2)(PERCISION) & MULTS_1_12_1(4,2)(PERCISION downto 1));
			MULTS_2_13_1(4,2)<=signed(MULTS_1_13_1(4,2)(PERCISION) & MULTS_1_13_1(4,2)(PERCISION downto 1));
			MULTS_2_14_1(4,2)<=signed(MULTS_1_14_1(4,2)(PERCISION) & MULTS_1_14_1(4,2)(PERCISION downto 1));
			MULTS_2_15_1(4,2)<=signed(MULTS_1_15_1(4,2)(PERCISION) & MULTS_1_15_1(4,2)(PERCISION downto 1));
			MULTS_2_16_1(4,2)<=signed(MULTS_1_16_1(4,2)(PERCISION) & MULTS_1_16_1(4,2)(PERCISION downto 1));

			MULTS_2_1_1(4,3)<=signed(MULTS_1_1_1(4,3)(PERCISION) & MULTS_1_1_1(4,3)(PERCISION downto 1));
			MULTS_2_2_1(4,3)<=signed(MULTS_1_2_1(4,3)(PERCISION) & MULTS_1_2_1(4,3)(PERCISION downto 1));
			MULTS_2_3_1(4,3)<=signed(MULTS_1_3_1(4,3)(PERCISION) & MULTS_1_3_1(4,3)(PERCISION downto 1));
			MULTS_2_4_1(4,3)<=signed(MULTS_1_4_1(4,3)(PERCISION) & MULTS_1_4_1(4,3)(PERCISION downto 1));
			MULTS_2_5_1(4,3)<=signed(MULTS_1_5_1(4,3)(PERCISION) & MULTS_1_5_1(4,3)(PERCISION downto 1));
			MULTS_2_6_1(4,3)<=signed(MULTS_1_6_1(4,3)(PERCISION) & MULTS_1_6_1(4,3)(PERCISION downto 1));
			MULTS_2_7_1(4,3)<=signed(MULTS_1_7_1(4,3)(PERCISION) & MULTS_1_7_1(4,3)(PERCISION downto 1));
			MULTS_2_8_1(4,3)<=signed(MULTS_1_8_1(4,3)(PERCISION) & MULTS_1_8_1(4,3)(PERCISION downto 1));
			MULTS_2_9_1(4,3)<=signed(MULTS_1_9_1(4,3)(PERCISION) & MULTS_1_9_1(4,3)(PERCISION downto 1));
			MULTS_2_10_1(4,3)<=signed(MULTS_1_10_1(4,3)(PERCISION) & MULTS_1_10_1(4,3)(PERCISION downto 1));
			MULTS_2_11_1(4,3)<=signed(MULTS_1_11_1(4,3)(PERCISION) & MULTS_1_11_1(4,3)(PERCISION downto 1));
			MULTS_2_12_1(4,3)<=signed(MULTS_1_12_1(4,3)(PERCISION) & MULTS_1_12_1(4,3)(PERCISION downto 1));
			MULTS_2_13_1(4,3)<=signed(MULTS_1_13_1(4,3)(PERCISION) & MULTS_1_13_1(4,3)(PERCISION downto 1));
			MULTS_2_14_1(4,3)<=signed(MULTS_1_14_1(4,3)(PERCISION) & MULTS_1_14_1(4,3)(PERCISION downto 1));
			MULTS_2_15_1(4,3)<=signed(MULTS_1_15_1(4,3)(PERCISION) & MULTS_1_15_1(4,3)(PERCISION downto 1));
			MULTS_2_16_1(4,3)<=signed(MULTS_1_16_1(4,3)(PERCISION) & MULTS_1_16_1(4,3)(PERCISION downto 1));

			MULTS_2_1_1(4,4)<=signed(MULTS_1_1_1(4,4)(PERCISION) & MULTS_1_1_1(4,4)(PERCISION downto 1));
			MULTS_2_2_1(4,4)<=signed(MULTS_1_2_1(4,4)(PERCISION) & MULTS_1_2_1(4,4)(PERCISION downto 1));
			MULTS_2_3_1(4,4)<=signed(MULTS_1_3_1(4,4)(PERCISION) & MULTS_1_3_1(4,4)(PERCISION downto 1));
			MULTS_2_4_1(4,4)<=signed(MULTS_1_4_1(4,4)(PERCISION) & MULTS_1_4_1(4,4)(PERCISION downto 1));
			MULTS_2_5_1(4,4)<=signed(MULTS_1_5_1(4,4)(PERCISION) & MULTS_1_5_1(4,4)(PERCISION downto 1));
			MULTS_2_6_1(4,4)<=signed(MULTS_1_6_1(4,4)(PERCISION) & MULTS_1_6_1(4,4)(PERCISION downto 1));
			MULTS_2_7_1(4,4)<=signed(MULTS_1_7_1(4,4)(PERCISION) & MULTS_1_7_1(4,4)(PERCISION downto 1));
			MULTS_2_8_1(4,4)<=signed(MULTS_1_8_1(4,4)(PERCISION) & MULTS_1_8_1(4,4)(PERCISION downto 1));
			MULTS_2_9_1(4,4)<=signed(MULTS_1_9_1(4,4)(PERCISION) & MULTS_1_9_1(4,4)(PERCISION downto 1));
			MULTS_2_10_1(4,4)<=signed(MULTS_1_10_1(4,4)(PERCISION) & MULTS_1_10_1(4,4)(PERCISION downto 1));
			MULTS_2_11_1(4,4)<=signed(MULTS_1_11_1(4,4)(PERCISION) & MULTS_1_11_1(4,4)(PERCISION downto 1));
			MULTS_2_12_1(4,4)<=signed(MULTS_1_12_1(4,4)(PERCISION) & MULTS_1_12_1(4,4)(PERCISION downto 1));
			MULTS_2_13_1(4,4)<=signed(MULTS_1_13_1(4,4)(PERCISION) & MULTS_1_13_1(4,4)(PERCISION downto 1));
			MULTS_2_14_1(4,4)<=signed(MULTS_1_14_1(4,4)(PERCISION) & MULTS_1_14_1(4,4)(PERCISION downto 1));
			MULTS_2_15_1(4,4)<=signed(MULTS_1_15_1(4,4)(PERCISION) & MULTS_1_15_1(4,4)(PERCISION downto 1));
			MULTS_2_16_1(4,4)<=signed(MULTS_1_16_1(4,4)(PERCISION) & MULTS_1_16_1(4,4)(PERCISION downto 1));

			MULTS_2_1_2(0,0)<=signed(MULTS_1_1_2(0,0)(PERCISION) & MULTS_1_1_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_1_3(0,0)(PERCISION) & MULTS_1_1_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(0,0)<=signed(MULTS_1_2_2(0,0)(PERCISION) & MULTS_1_2_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_2_3(0,0)(PERCISION) & MULTS_1_2_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(0,0)<=signed(MULTS_1_3_2(0,0)(PERCISION) & MULTS_1_3_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_3_3(0,0)(PERCISION) & MULTS_1_3_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(0,0)<=signed(MULTS_1_4_2(0,0)(PERCISION) & MULTS_1_4_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_4_3(0,0)(PERCISION) & MULTS_1_4_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(0,0)<=signed(MULTS_1_5_2(0,0)(PERCISION) & MULTS_1_5_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_5_3(0,0)(PERCISION) & MULTS_1_5_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(0,0)<=signed(MULTS_1_6_2(0,0)(PERCISION) & MULTS_1_6_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_6_3(0,0)(PERCISION) & MULTS_1_6_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(0,0)<=signed(MULTS_1_7_2(0,0)(PERCISION) & MULTS_1_7_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_7_3(0,0)(PERCISION) & MULTS_1_7_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(0,0)<=signed(MULTS_1_8_2(0,0)(PERCISION) & MULTS_1_8_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_8_3(0,0)(PERCISION) & MULTS_1_8_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(0,0)<=signed(MULTS_1_9_2(0,0)(PERCISION) & MULTS_1_9_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_9_3(0,0)(PERCISION) & MULTS_1_9_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(0,0)<=signed(MULTS_1_10_2(0,0)(PERCISION) & MULTS_1_10_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_10_3(0,0)(PERCISION) & MULTS_1_10_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(0,0)<=signed(MULTS_1_11_2(0,0)(PERCISION) & MULTS_1_11_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_11_3(0,0)(PERCISION) & MULTS_1_11_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(0,0)<=signed(MULTS_1_12_2(0,0)(PERCISION) & MULTS_1_12_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_12_3(0,0)(PERCISION) & MULTS_1_12_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(0,0)<=signed(MULTS_1_13_2(0,0)(PERCISION) & MULTS_1_13_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_13_3(0,0)(PERCISION) & MULTS_1_13_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(0,0)<=signed(MULTS_1_14_2(0,0)(PERCISION) & MULTS_1_14_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_14_3(0,0)(PERCISION) & MULTS_1_14_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(0,0)<=signed(MULTS_1_15_2(0,0)(PERCISION) & MULTS_1_15_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_15_3(0,0)(PERCISION) & MULTS_1_15_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(0,0)<=signed(MULTS_1_16_2(0,0)(PERCISION) & MULTS_1_16_2(0,0)(PERCISION downto 1)) + signed(MULTS_1_16_3(0,0)(PERCISION) & MULTS_1_16_3(0,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(0,0) ------------------

			MULTS_2_1_2(0,1)<=signed(MULTS_1_1_2(0,1)(PERCISION) & MULTS_1_1_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_1_3(0,1)(PERCISION) & MULTS_1_1_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(0,1)<=signed(MULTS_1_2_2(0,1)(PERCISION) & MULTS_1_2_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_2_3(0,1)(PERCISION) & MULTS_1_2_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(0,1)<=signed(MULTS_1_3_2(0,1)(PERCISION) & MULTS_1_3_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_3_3(0,1)(PERCISION) & MULTS_1_3_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(0,1)<=signed(MULTS_1_4_2(0,1)(PERCISION) & MULTS_1_4_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_4_3(0,1)(PERCISION) & MULTS_1_4_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(0,1)<=signed(MULTS_1_5_2(0,1)(PERCISION) & MULTS_1_5_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_5_3(0,1)(PERCISION) & MULTS_1_5_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(0,1)<=signed(MULTS_1_6_2(0,1)(PERCISION) & MULTS_1_6_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_6_3(0,1)(PERCISION) & MULTS_1_6_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(0,1)<=signed(MULTS_1_7_2(0,1)(PERCISION) & MULTS_1_7_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_7_3(0,1)(PERCISION) & MULTS_1_7_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(0,1)<=signed(MULTS_1_8_2(0,1)(PERCISION) & MULTS_1_8_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_8_3(0,1)(PERCISION) & MULTS_1_8_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(0,1)<=signed(MULTS_1_9_2(0,1)(PERCISION) & MULTS_1_9_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_9_3(0,1)(PERCISION) & MULTS_1_9_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(0,1)<=signed(MULTS_1_10_2(0,1)(PERCISION) & MULTS_1_10_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_10_3(0,1)(PERCISION) & MULTS_1_10_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(0,1)<=signed(MULTS_1_11_2(0,1)(PERCISION) & MULTS_1_11_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_11_3(0,1)(PERCISION) & MULTS_1_11_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(0,1)<=signed(MULTS_1_12_2(0,1)(PERCISION) & MULTS_1_12_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_12_3(0,1)(PERCISION) & MULTS_1_12_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(0,1)<=signed(MULTS_1_13_2(0,1)(PERCISION) & MULTS_1_13_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_13_3(0,1)(PERCISION) & MULTS_1_13_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(0,1)<=signed(MULTS_1_14_2(0,1)(PERCISION) & MULTS_1_14_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_14_3(0,1)(PERCISION) & MULTS_1_14_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(0,1)<=signed(MULTS_1_15_2(0,1)(PERCISION) & MULTS_1_15_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_15_3(0,1)(PERCISION) & MULTS_1_15_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(0,1)<=signed(MULTS_1_16_2(0,1)(PERCISION) & MULTS_1_16_2(0,1)(PERCISION downto 1)) + signed(MULTS_1_16_3(0,1)(PERCISION) & MULTS_1_16_3(0,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(0,1) ------------------

			MULTS_2_1_2(0,2)<=signed(MULTS_1_1_2(0,2)(PERCISION) & MULTS_1_1_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_1_3(0,2)(PERCISION) & MULTS_1_1_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(0,2)<=signed(MULTS_1_2_2(0,2)(PERCISION) & MULTS_1_2_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_2_3(0,2)(PERCISION) & MULTS_1_2_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(0,2)<=signed(MULTS_1_3_2(0,2)(PERCISION) & MULTS_1_3_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_3_3(0,2)(PERCISION) & MULTS_1_3_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(0,2)<=signed(MULTS_1_4_2(0,2)(PERCISION) & MULTS_1_4_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_4_3(0,2)(PERCISION) & MULTS_1_4_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(0,2)<=signed(MULTS_1_5_2(0,2)(PERCISION) & MULTS_1_5_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_5_3(0,2)(PERCISION) & MULTS_1_5_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(0,2)<=signed(MULTS_1_6_2(0,2)(PERCISION) & MULTS_1_6_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_6_3(0,2)(PERCISION) & MULTS_1_6_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(0,2)<=signed(MULTS_1_7_2(0,2)(PERCISION) & MULTS_1_7_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_7_3(0,2)(PERCISION) & MULTS_1_7_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(0,2)<=signed(MULTS_1_8_2(0,2)(PERCISION) & MULTS_1_8_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_8_3(0,2)(PERCISION) & MULTS_1_8_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(0,2)<=signed(MULTS_1_9_2(0,2)(PERCISION) & MULTS_1_9_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_9_3(0,2)(PERCISION) & MULTS_1_9_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(0,2)<=signed(MULTS_1_10_2(0,2)(PERCISION) & MULTS_1_10_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_10_3(0,2)(PERCISION) & MULTS_1_10_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(0,2)<=signed(MULTS_1_11_2(0,2)(PERCISION) & MULTS_1_11_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_11_3(0,2)(PERCISION) & MULTS_1_11_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(0,2)<=signed(MULTS_1_12_2(0,2)(PERCISION) & MULTS_1_12_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_12_3(0,2)(PERCISION) & MULTS_1_12_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(0,2)<=signed(MULTS_1_13_2(0,2)(PERCISION) & MULTS_1_13_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_13_3(0,2)(PERCISION) & MULTS_1_13_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(0,2)<=signed(MULTS_1_14_2(0,2)(PERCISION) & MULTS_1_14_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_14_3(0,2)(PERCISION) & MULTS_1_14_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(0,2)<=signed(MULTS_1_15_2(0,2)(PERCISION) & MULTS_1_15_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_15_3(0,2)(PERCISION) & MULTS_1_15_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(0,2)<=signed(MULTS_1_16_2(0,2)(PERCISION) & MULTS_1_16_2(0,2)(PERCISION downto 1)) + signed(MULTS_1_16_3(0,2)(PERCISION) & MULTS_1_16_3(0,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(0,2) ------------------

			MULTS_2_1_2(0,3)<=signed(MULTS_1_1_2(0,3)(PERCISION) & MULTS_1_1_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_1_3(0,3)(PERCISION) & MULTS_1_1_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(0,3)<=signed(MULTS_1_2_2(0,3)(PERCISION) & MULTS_1_2_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_2_3(0,3)(PERCISION) & MULTS_1_2_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(0,3)<=signed(MULTS_1_3_2(0,3)(PERCISION) & MULTS_1_3_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_3_3(0,3)(PERCISION) & MULTS_1_3_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(0,3)<=signed(MULTS_1_4_2(0,3)(PERCISION) & MULTS_1_4_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_4_3(0,3)(PERCISION) & MULTS_1_4_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(0,3)<=signed(MULTS_1_5_2(0,3)(PERCISION) & MULTS_1_5_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_5_3(0,3)(PERCISION) & MULTS_1_5_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(0,3)<=signed(MULTS_1_6_2(0,3)(PERCISION) & MULTS_1_6_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_6_3(0,3)(PERCISION) & MULTS_1_6_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(0,3)<=signed(MULTS_1_7_2(0,3)(PERCISION) & MULTS_1_7_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_7_3(0,3)(PERCISION) & MULTS_1_7_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(0,3)<=signed(MULTS_1_8_2(0,3)(PERCISION) & MULTS_1_8_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_8_3(0,3)(PERCISION) & MULTS_1_8_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(0,3)<=signed(MULTS_1_9_2(0,3)(PERCISION) & MULTS_1_9_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_9_3(0,3)(PERCISION) & MULTS_1_9_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(0,3)<=signed(MULTS_1_10_2(0,3)(PERCISION) & MULTS_1_10_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_10_3(0,3)(PERCISION) & MULTS_1_10_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(0,3)<=signed(MULTS_1_11_2(0,3)(PERCISION) & MULTS_1_11_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_11_3(0,3)(PERCISION) & MULTS_1_11_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(0,3)<=signed(MULTS_1_12_2(0,3)(PERCISION) & MULTS_1_12_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_12_3(0,3)(PERCISION) & MULTS_1_12_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(0,3)<=signed(MULTS_1_13_2(0,3)(PERCISION) & MULTS_1_13_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_13_3(0,3)(PERCISION) & MULTS_1_13_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(0,3)<=signed(MULTS_1_14_2(0,3)(PERCISION) & MULTS_1_14_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_14_3(0,3)(PERCISION) & MULTS_1_14_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(0,3)<=signed(MULTS_1_15_2(0,3)(PERCISION) & MULTS_1_15_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_15_3(0,3)(PERCISION) & MULTS_1_15_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(0,3)<=signed(MULTS_1_16_2(0,3)(PERCISION) & MULTS_1_16_2(0,3)(PERCISION downto 1)) + signed(MULTS_1_16_3(0,3)(PERCISION) & MULTS_1_16_3(0,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(0,3) ------------------

			MULTS_2_1_2(0,4)<=signed(MULTS_1_1_2(0,4)(PERCISION) & MULTS_1_1_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_1_3(0,4)(PERCISION) & MULTS_1_1_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(0,4)<=signed(MULTS_1_2_2(0,4)(PERCISION) & MULTS_1_2_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_2_3(0,4)(PERCISION) & MULTS_1_2_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(0,4)<=signed(MULTS_1_3_2(0,4)(PERCISION) & MULTS_1_3_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_3_3(0,4)(PERCISION) & MULTS_1_3_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(0,4)<=signed(MULTS_1_4_2(0,4)(PERCISION) & MULTS_1_4_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_4_3(0,4)(PERCISION) & MULTS_1_4_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(0,4)<=signed(MULTS_1_5_2(0,4)(PERCISION) & MULTS_1_5_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_5_3(0,4)(PERCISION) & MULTS_1_5_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(0,4)<=signed(MULTS_1_6_2(0,4)(PERCISION) & MULTS_1_6_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_6_3(0,4)(PERCISION) & MULTS_1_6_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(0,4)<=signed(MULTS_1_7_2(0,4)(PERCISION) & MULTS_1_7_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_7_3(0,4)(PERCISION) & MULTS_1_7_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(0,4)<=signed(MULTS_1_8_2(0,4)(PERCISION) & MULTS_1_8_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_8_3(0,4)(PERCISION) & MULTS_1_8_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(0,4)<=signed(MULTS_1_9_2(0,4)(PERCISION) & MULTS_1_9_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_9_3(0,4)(PERCISION) & MULTS_1_9_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(0,4)<=signed(MULTS_1_10_2(0,4)(PERCISION) & MULTS_1_10_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_10_3(0,4)(PERCISION) & MULTS_1_10_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(0,4)<=signed(MULTS_1_11_2(0,4)(PERCISION) & MULTS_1_11_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_11_3(0,4)(PERCISION) & MULTS_1_11_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(0,4)<=signed(MULTS_1_12_2(0,4)(PERCISION) & MULTS_1_12_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_12_3(0,4)(PERCISION) & MULTS_1_12_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(0,4)<=signed(MULTS_1_13_2(0,4)(PERCISION) & MULTS_1_13_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_13_3(0,4)(PERCISION) & MULTS_1_13_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(0,4)<=signed(MULTS_1_14_2(0,4)(PERCISION) & MULTS_1_14_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_14_3(0,4)(PERCISION) & MULTS_1_14_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(0,4)<=signed(MULTS_1_15_2(0,4)(PERCISION) & MULTS_1_15_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_15_3(0,4)(PERCISION) & MULTS_1_15_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(0,4)<=signed(MULTS_1_16_2(0,4)(PERCISION) & MULTS_1_16_2(0,4)(PERCISION downto 1)) + signed(MULTS_1_16_3(0,4)(PERCISION) & MULTS_1_16_3(0,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(0,4) ------------------

			MULTS_2_1_2(1,0)<=signed(MULTS_1_1_2(1,0)(PERCISION) & MULTS_1_1_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_1_3(1,0)(PERCISION) & MULTS_1_1_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(1,0)<=signed(MULTS_1_2_2(1,0)(PERCISION) & MULTS_1_2_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_2_3(1,0)(PERCISION) & MULTS_1_2_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(1,0)<=signed(MULTS_1_3_2(1,0)(PERCISION) & MULTS_1_3_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_3_3(1,0)(PERCISION) & MULTS_1_3_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(1,0)<=signed(MULTS_1_4_2(1,0)(PERCISION) & MULTS_1_4_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_4_3(1,0)(PERCISION) & MULTS_1_4_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(1,0)<=signed(MULTS_1_5_2(1,0)(PERCISION) & MULTS_1_5_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_5_3(1,0)(PERCISION) & MULTS_1_5_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(1,0)<=signed(MULTS_1_6_2(1,0)(PERCISION) & MULTS_1_6_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_6_3(1,0)(PERCISION) & MULTS_1_6_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(1,0)<=signed(MULTS_1_7_2(1,0)(PERCISION) & MULTS_1_7_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_7_3(1,0)(PERCISION) & MULTS_1_7_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(1,0)<=signed(MULTS_1_8_2(1,0)(PERCISION) & MULTS_1_8_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_8_3(1,0)(PERCISION) & MULTS_1_8_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(1,0)<=signed(MULTS_1_9_2(1,0)(PERCISION) & MULTS_1_9_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_9_3(1,0)(PERCISION) & MULTS_1_9_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(1,0)<=signed(MULTS_1_10_2(1,0)(PERCISION) & MULTS_1_10_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_10_3(1,0)(PERCISION) & MULTS_1_10_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(1,0)<=signed(MULTS_1_11_2(1,0)(PERCISION) & MULTS_1_11_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_11_3(1,0)(PERCISION) & MULTS_1_11_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(1,0)<=signed(MULTS_1_12_2(1,0)(PERCISION) & MULTS_1_12_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_12_3(1,0)(PERCISION) & MULTS_1_12_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(1,0)<=signed(MULTS_1_13_2(1,0)(PERCISION) & MULTS_1_13_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_13_3(1,0)(PERCISION) & MULTS_1_13_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(1,0)<=signed(MULTS_1_14_2(1,0)(PERCISION) & MULTS_1_14_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_14_3(1,0)(PERCISION) & MULTS_1_14_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(1,0)<=signed(MULTS_1_15_2(1,0)(PERCISION) & MULTS_1_15_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_15_3(1,0)(PERCISION) & MULTS_1_15_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(1,0)<=signed(MULTS_1_16_2(1,0)(PERCISION) & MULTS_1_16_2(1,0)(PERCISION downto 1)) + signed(MULTS_1_16_3(1,0)(PERCISION) & MULTS_1_16_3(1,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(1,0) ------------------

			MULTS_2_1_2(1,1)<=signed(MULTS_1_1_2(1,1)(PERCISION) & MULTS_1_1_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_1_3(1,1)(PERCISION) & MULTS_1_1_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(1,1)<=signed(MULTS_1_2_2(1,1)(PERCISION) & MULTS_1_2_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_2_3(1,1)(PERCISION) & MULTS_1_2_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(1,1)<=signed(MULTS_1_3_2(1,1)(PERCISION) & MULTS_1_3_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_3_3(1,1)(PERCISION) & MULTS_1_3_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(1,1)<=signed(MULTS_1_4_2(1,1)(PERCISION) & MULTS_1_4_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_4_3(1,1)(PERCISION) & MULTS_1_4_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(1,1)<=signed(MULTS_1_5_2(1,1)(PERCISION) & MULTS_1_5_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_5_3(1,1)(PERCISION) & MULTS_1_5_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(1,1)<=signed(MULTS_1_6_2(1,1)(PERCISION) & MULTS_1_6_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_6_3(1,1)(PERCISION) & MULTS_1_6_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(1,1)<=signed(MULTS_1_7_2(1,1)(PERCISION) & MULTS_1_7_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_7_3(1,1)(PERCISION) & MULTS_1_7_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(1,1)<=signed(MULTS_1_8_2(1,1)(PERCISION) & MULTS_1_8_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_8_3(1,1)(PERCISION) & MULTS_1_8_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(1,1)<=signed(MULTS_1_9_2(1,1)(PERCISION) & MULTS_1_9_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_9_3(1,1)(PERCISION) & MULTS_1_9_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(1,1)<=signed(MULTS_1_10_2(1,1)(PERCISION) & MULTS_1_10_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_10_3(1,1)(PERCISION) & MULTS_1_10_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(1,1)<=signed(MULTS_1_11_2(1,1)(PERCISION) & MULTS_1_11_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_11_3(1,1)(PERCISION) & MULTS_1_11_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(1,1)<=signed(MULTS_1_12_2(1,1)(PERCISION) & MULTS_1_12_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_12_3(1,1)(PERCISION) & MULTS_1_12_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(1,1)<=signed(MULTS_1_13_2(1,1)(PERCISION) & MULTS_1_13_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_13_3(1,1)(PERCISION) & MULTS_1_13_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(1,1)<=signed(MULTS_1_14_2(1,1)(PERCISION) & MULTS_1_14_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_14_3(1,1)(PERCISION) & MULTS_1_14_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(1,1)<=signed(MULTS_1_15_2(1,1)(PERCISION) & MULTS_1_15_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_15_3(1,1)(PERCISION) & MULTS_1_15_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(1,1)<=signed(MULTS_1_16_2(1,1)(PERCISION) & MULTS_1_16_2(1,1)(PERCISION downto 1)) + signed(MULTS_1_16_3(1,1)(PERCISION) & MULTS_1_16_3(1,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(1,1) ------------------

			MULTS_2_1_2(1,2)<=signed(MULTS_1_1_2(1,2)(PERCISION) & MULTS_1_1_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_1_3(1,2)(PERCISION) & MULTS_1_1_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(1,2)<=signed(MULTS_1_2_2(1,2)(PERCISION) & MULTS_1_2_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_2_3(1,2)(PERCISION) & MULTS_1_2_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(1,2)<=signed(MULTS_1_3_2(1,2)(PERCISION) & MULTS_1_3_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_3_3(1,2)(PERCISION) & MULTS_1_3_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(1,2)<=signed(MULTS_1_4_2(1,2)(PERCISION) & MULTS_1_4_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_4_3(1,2)(PERCISION) & MULTS_1_4_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(1,2)<=signed(MULTS_1_5_2(1,2)(PERCISION) & MULTS_1_5_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_5_3(1,2)(PERCISION) & MULTS_1_5_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(1,2)<=signed(MULTS_1_6_2(1,2)(PERCISION) & MULTS_1_6_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_6_3(1,2)(PERCISION) & MULTS_1_6_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(1,2)<=signed(MULTS_1_7_2(1,2)(PERCISION) & MULTS_1_7_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_7_3(1,2)(PERCISION) & MULTS_1_7_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(1,2)<=signed(MULTS_1_8_2(1,2)(PERCISION) & MULTS_1_8_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_8_3(1,2)(PERCISION) & MULTS_1_8_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(1,2)<=signed(MULTS_1_9_2(1,2)(PERCISION) & MULTS_1_9_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_9_3(1,2)(PERCISION) & MULTS_1_9_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(1,2)<=signed(MULTS_1_10_2(1,2)(PERCISION) & MULTS_1_10_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_10_3(1,2)(PERCISION) & MULTS_1_10_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(1,2)<=signed(MULTS_1_11_2(1,2)(PERCISION) & MULTS_1_11_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_11_3(1,2)(PERCISION) & MULTS_1_11_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(1,2)<=signed(MULTS_1_12_2(1,2)(PERCISION) & MULTS_1_12_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_12_3(1,2)(PERCISION) & MULTS_1_12_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(1,2)<=signed(MULTS_1_13_2(1,2)(PERCISION) & MULTS_1_13_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_13_3(1,2)(PERCISION) & MULTS_1_13_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(1,2)<=signed(MULTS_1_14_2(1,2)(PERCISION) & MULTS_1_14_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_14_3(1,2)(PERCISION) & MULTS_1_14_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(1,2)<=signed(MULTS_1_15_2(1,2)(PERCISION) & MULTS_1_15_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_15_3(1,2)(PERCISION) & MULTS_1_15_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(1,2)<=signed(MULTS_1_16_2(1,2)(PERCISION) & MULTS_1_16_2(1,2)(PERCISION downto 1)) + signed(MULTS_1_16_3(1,2)(PERCISION) & MULTS_1_16_3(1,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(1,2) ------------------

			MULTS_2_1_2(1,3)<=signed(MULTS_1_1_2(1,3)(PERCISION) & MULTS_1_1_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_1_3(1,3)(PERCISION) & MULTS_1_1_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(1,3)<=signed(MULTS_1_2_2(1,3)(PERCISION) & MULTS_1_2_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_2_3(1,3)(PERCISION) & MULTS_1_2_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(1,3)<=signed(MULTS_1_3_2(1,3)(PERCISION) & MULTS_1_3_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_3_3(1,3)(PERCISION) & MULTS_1_3_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(1,3)<=signed(MULTS_1_4_2(1,3)(PERCISION) & MULTS_1_4_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_4_3(1,3)(PERCISION) & MULTS_1_4_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(1,3)<=signed(MULTS_1_5_2(1,3)(PERCISION) & MULTS_1_5_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_5_3(1,3)(PERCISION) & MULTS_1_5_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(1,3)<=signed(MULTS_1_6_2(1,3)(PERCISION) & MULTS_1_6_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_6_3(1,3)(PERCISION) & MULTS_1_6_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(1,3)<=signed(MULTS_1_7_2(1,3)(PERCISION) & MULTS_1_7_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_7_3(1,3)(PERCISION) & MULTS_1_7_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(1,3)<=signed(MULTS_1_8_2(1,3)(PERCISION) & MULTS_1_8_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_8_3(1,3)(PERCISION) & MULTS_1_8_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(1,3)<=signed(MULTS_1_9_2(1,3)(PERCISION) & MULTS_1_9_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_9_3(1,3)(PERCISION) & MULTS_1_9_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(1,3)<=signed(MULTS_1_10_2(1,3)(PERCISION) & MULTS_1_10_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_10_3(1,3)(PERCISION) & MULTS_1_10_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(1,3)<=signed(MULTS_1_11_2(1,3)(PERCISION) & MULTS_1_11_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_11_3(1,3)(PERCISION) & MULTS_1_11_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(1,3)<=signed(MULTS_1_12_2(1,3)(PERCISION) & MULTS_1_12_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_12_3(1,3)(PERCISION) & MULTS_1_12_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(1,3)<=signed(MULTS_1_13_2(1,3)(PERCISION) & MULTS_1_13_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_13_3(1,3)(PERCISION) & MULTS_1_13_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(1,3)<=signed(MULTS_1_14_2(1,3)(PERCISION) & MULTS_1_14_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_14_3(1,3)(PERCISION) & MULTS_1_14_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(1,3)<=signed(MULTS_1_15_2(1,3)(PERCISION) & MULTS_1_15_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_15_3(1,3)(PERCISION) & MULTS_1_15_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(1,3)<=signed(MULTS_1_16_2(1,3)(PERCISION) & MULTS_1_16_2(1,3)(PERCISION downto 1)) + signed(MULTS_1_16_3(1,3)(PERCISION) & MULTS_1_16_3(1,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(1,3) ------------------

			MULTS_2_1_2(1,4)<=signed(MULTS_1_1_2(1,4)(PERCISION) & MULTS_1_1_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_1_3(1,4)(PERCISION) & MULTS_1_1_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(1,4)<=signed(MULTS_1_2_2(1,4)(PERCISION) & MULTS_1_2_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_2_3(1,4)(PERCISION) & MULTS_1_2_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(1,4)<=signed(MULTS_1_3_2(1,4)(PERCISION) & MULTS_1_3_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_3_3(1,4)(PERCISION) & MULTS_1_3_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(1,4)<=signed(MULTS_1_4_2(1,4)(PERCISION) & MULTS_1_4_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_4_3(1,4)(PERCISION) & MULTS_1_4_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(1,4)<=signed(MULTS_1_5_2(1,4)(PERCISION) & MULTS_1_5_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_5_3(1,4)(PERCISION) & MULTS_1_5_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(1,4)<=signed(MULTS_1_6_2(1,4)(PERCISION) & MULTS_1_6_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_6_3(1,4)(PERCISION) & MULTS_1_6_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(1,4)<=signed(MULTS_1_7_2(1,4)(PERCISION) & MULTS_1_7_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_7_3(1,4)(PERCISION) & MULTS_1_7_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(1,4)<=signed(MULTS_1_8_2(1,4)(PERCISION) & MULTS_1_8_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_8_3(1,4)(PERCISION) & MULTS_1_8_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(1,4)<=signed(MULTS_1_9_2(1,4)(PERCISION) & MULTS_1_9_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_9_3(1,4)(PERCISION) & MULTS_1_9_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(1,4)<=signed(MULTS_1_10_2(1,4)(PERCISION) & MULTS_1_10_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_10_3(1,4)(PERCISION) & MULTS_1_10_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(1,4)<=signed(MULTS_1_11_2(1,4)(PERCISION) & MULTS_1_11_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_11_3(1,4)(PERCISION) & MULTS_1_11_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(1,4)<=signed(MULTS_1_12_2(1,4)(PERCISION) & MULTS_1_12_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_12_3(1,4)(PERCISION) & MULTS_1_12_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(1,4)<=signed(MULTS_1_13_2(1,4)(PERCISION) & MULTS_1_13_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_13_3(1,4)(PERCISION) & MULTS_1_13_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(1,4)<=signed(MULTS_1_14_2(1,4)(PERCISION) & MULTS_1_14_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_14_3(1,4)(PERCISION) & MULTS_1_14_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(1,4)<=signed(MULTS_1_15_2(1,4)(PERCISION) & MULTS_1_15_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_15_3(1,4)(PERCISION) & MULTS_1_15_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(1,4)<=signed(MULTS_1_16_2(1,4)(PERCISION) & MULTS_1_16_2(1,4)(PERCISION downto 1)) + signed(MULTS_1_16_3(1,4)(PERCISION) & MULTS_1_16_3(1,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(1,4) ------------------

			MULTS_2_1_2(2,0)<=signed(MULTS_1_1_2(2,0)(PERCISION) & MULTS_1_1_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_1_3(2,0)(PERCISION) & MULTS_1_1_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(2,0)<=signed(MULTS_1_2_2(2,0)(PERCISION) & MULTS_1_2_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_2_3(2,0)(PERCISION) & MULTS_1_2_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(2,0)<=signed(MULTS_1_3_2(2,0)(PERCISION) & MULTS_1_3_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_3_3(2,0)(PERCISION) & MULTS_1_3_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(2,0)<=signed(MULTS_1_4_2(2,0)(PERCISION) & MULTS_1_4_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_4_3(2,0)(PERCISION) & MULTS_1_4_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(2,0)<=signed(MULTS_1_5_2(2,0)(PERCISION) & MULTS_1_5_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_5_3(2,0)(PERCISION) & MULTS_1_5_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(2,0)<=signed(MULTS_1_6_2(2,0)(PERCISION) & MULTS_1_6_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_6_3(2,0)(PERCISION) & MULTS_1_6_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(2,0)<=signed(MULTS_1_7_2(2,0)(PERCISION) & MULTS_1_7_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_7_3(2,0)(PERCISION) & MULTS_1_7_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(2,0)<=signed(MULTS_1_8_2(2,0)(PERCISION) & MULTS_1_8_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_8_3(2,0)(PERCISION) & MULTS_1_8_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(2,0)<=signed(MULTS_1_9_2(2,0)(PERCISION) & MULTS_1_9_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_9_3(2,0)(PERCISION) & MULTS_1_9_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(2,0)<=signed(MULTS_1_10_2(2,0)(PERCISION) & MULTS_1_10_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_10_3(2,0)(PERCISION) & MULTS_1_10_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(2,0)<=signed(MULTS_1_11_2(2,0)(PERCISION) & MULTS_1_11_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_11_3(2,0)(PERCISION) & MULTS_1_11_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(2,0)<=signed(MULTS_1_12_2(2,0)(PERCISION) & MULTS_1_12_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_12_3(2,0)(PERCISION) & MULTS_1_12_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(2,0)<=signed(MULTS_1_13_2(2,0)(PERCISION) & MULTS_1_13_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_13_3(2,0)(PERCISION) & MULTS_1_13_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(2,0)<=signed(MULTS_1_14_2(2,0)(PERCISION) & MULTS_1_14_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_14_3(2,0)(PERCISION) & MULTS_1_14_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(2,0)<=signed(MULTS_1_15_2(2,0)(PERCISION) & MULTS_1_15_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_15_3(2,0)(PERCISION) & MULTS_1_15_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(2,0)<=signed(MULTS_1_16_2(2,0)(PERCISION) & MULTS_1_16_2(2,0)(PERCISION downto 1)) + signed(MULTS_1_16_3(2,0)(PERCISION) & MULTS_1_16_3(2,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(2,0) ------------------

			MULTS_2_1_2(2,1)<=signed(MULTS_1_1_2(2,1)(PERCISION) & MULTS_1_1_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_1_3(2,1)(PERCISION) & MULTS_1_1_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(2,1)<=signed(MULTS_1_2_2(2,1)(PERCISION) & MULTS_1_2_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_2_3(2,1)(PERCISION) & MULTS_1_2_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(2,1)<=signed(MULTS_1_3_2(2,1)(PERCISION) & MULTS_1_3_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_3_3(2,1)(PERCISION) & MULTS_1_3_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(2,1)<=signed(MULTS_1_4_2(2,1)(PERCISION) & MULTS_1_4_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_4_3(2,1)(PERCISION) & MULTS_1_4_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(2,1)<=signed(MULTS_1_5_2(2,1)(PERCISION) & MULTS_1_5_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_5_3(2,1)(PERCISION) & MULTS_1_5_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(2,1)<=signed(MULTS_1_6_2(2,1)(PERCISION) & MULTS_1_6_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_6_3(2,1)(PERCISION) & MULTS_1_6_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(2,1)<=signed(MULTS_1_7_2(2,1)(PERCISION) & MULTS_1_7_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_7_3(2,1)(PERCISION) & MULTS_1_7_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(2,1)<=signed(MULTS_1_8_2(2,1)(PERCISION) & MULTS_1_8_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_8_3(2,1)(PERCISION) & MULTS_1_8_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(2,1)<=signed(MULTS_1_9_2(2,1)(PERCISION) & MULTS_1_9_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_9_3(2,1)(PERCISION) & MULTS_1_9_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(2,1)<=signed(MULTS_1_10_2(2,1)(PERCISION) & MULTS_1_10_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_10_3(2,1)(PERCISION) & MULTS_1_10_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(2,1)<=signed(MULTS_1_11_2(2,1)(PERCISION) & MULTS_1_11_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_11_3(2,1)(PERCISION) & MULTS_1_11_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(2,1)<=signed(MULTS_1_12_2(2,1)(PERCISION) & MULTS_1_12_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_12_3(2,1)(PERCISION) & MULTS_1_12_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(2,1)<=signed(MULTS_1_13_2(2,1)(PERCISION) & MULTS_1_13_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_13_3(2,1)(PERCISION) & MULTS_1_13_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(2,1)<=signed(MULTS_1_14_2(2,1)(PERCISION) & MULTS_1_14_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_14_3(2,1)(PERCISION) & MULTS_1_14_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(2,1)<=signed(MULTS_1_15_2(2,1)(PERCISION) & MULTS_1_15_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_15_3(2,1)(PERCISION) & MULTS_1_15_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(2,1)<=signed(MULTS_1_16_2(2,1)(PERCISION) & MULTS_1_16_2(2,1)(PERCISION downto 1)) + signed(MULTS_1_16_3(2,1)(PERCISION) & MULTS_1_16_3(2,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(2,1) ------------------

			MULTS_2_1_2(2,2)<=signed(MULTS_1_1_2(2,2)(PERCISION) & MULTS_1_1_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_1_3(2,2)(PERCISION) & MULTS_1_1_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(2,2)<=signed(MULTS_1_2_2(2,2)(PERCISION) & MULTS_1_2_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_2_3(2,2)(PERCISION) & MULTS_1_2_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(2,2)<=signed(MULTS_1_3_2(2,2)(PERCISION) & MULTS_1_3_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_3_3(2,2)(PERCISION) & MULTS_1_3_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(2,2)<=signed(MULTS_1_4_2(2,2)(PERCISION) & MULTS_1_4_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_4_3(2,2)(PERCISION) & MULTS_1_4_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(2,2)<=signed(MULTS_1_5_2(2,2)(PERCISION) & MULTS_1_5_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_5_3(2,2)(PERCISION) & MULTS_1_5_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(2,2)<=signed(MULTS_1_6_2(2,2)(PERCISION) & MULTS_1_6_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_6_3(2,2)(PERCISION) & MULTS_1_6_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(2,2)<=signed(MULTS_1_7_2(2,2)(PERCISION) & MULTS_1_7_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_7_3(2,2)(PERCISION) & MULTS_1_7_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(2,2)<=signed(MULTS_1_8_2(2,2)(PERCISION) & MULTS_1_8_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_8_3(2,2)(PERCISION) & MULTS_1_8_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(2,2)<=signed(MULTS_1_9_2(2,2)(PERCISION) & MULTS_1_9_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_9_3(2,2)(PERCISION) & MULTS_1_9_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(2,2)<=signed(MULTS_1_10_2(2,2)(PERCISION) & MULTS_1_10_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_10_3(2,2)(PERCISION) & MULTS_1_10_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(2,2)<=signed(MULTS_1_11_2(2,2)(PERCISION) & MULTS_1_11_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_11_3(2,2)(PERCISION) & MULTS_1_11_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(2,2)<=signed(MULTS_1_12_2(2,2)(PERCISION) & MULTS_1_12_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_12_3(2,2)(PERCISION) & MULTS_1_12_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(2,2)<=signed(MULTS_1_13_2(2,2)(PERCISION) & MULTS_1_13_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_13_3(2,2)(PERCISION) & MULTS_1_13_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(2,2)<=signed(MULTS_1_14_2(2,2)(PERCISION) & MULTS_1_14_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_14_3(2,2)(PERCISION) & MULTS_1_14_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(2,2)<=signed(MULTS_1_15_2(2,2)(PERCISION) & MULTS_1_15_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_15_3(2,2)(PERCISION) & MULTS_1_15_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(2,2)<=signed(MULTS_1_16_2(2,2)(PERCISION) & MULTS_1_16_2(2,2)(PERCISION downto 1)) + signed(MULTS_1_16_3(2,2)(PERCISION) & MULTS_1_16_3(2,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(2,2) ------------------

			MULTS_2_1_2(2,3)<=signed(MULTS_1_1_2(2,3)(PERCISION) & MULTS_1_1_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_1_3(2,3)(PERCISION) & MULTS_1_1_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(2,3)<=signed(MULTS_1_2_2(2,3)(PERCISION) & MULTS_1_2_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_2_3(2,3)(PERCISION) & MULTS_1_2_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(2,3)<=signed(MULTS_1_3_2(2,3)(PERCISION) & MULTS_1_3_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_3_3(2,3)(PERCISION) & MULTS_1_3_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(2,3)<=signed(MULTS_1_4_2(2,3)(PERCISION) & MULTS_1_4_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_4_3(2,3)(PERCISION) & MULTS_1_4_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(2,3)<=signed(MULTS_1_5_2(2,3)(PERCISION) & MULTS_1_5_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_5_3(2,3)(PERCISION) & MULTS_1_5_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(2,3)<=signed(MULTS_1_6_2(2,3)(PERCISION) & MULTS_1_6_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_6_3(2,3)(PERCISION) & MULTS_1_6_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(2,3)<=signed(MULTS_1_7_2(2,3)(PERCISION) & MULTS_1_7_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_7_3(2,3)(PERCISION) & MULTS_1_7_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(2,3)<=signed(MULTS_1_8_2(2,3)(PERCISION) & MULTS_1_8_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_8_3(2,3)(PERCISION) & MULTS_1_8_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(2,3)<=signed(MULTS_1_9_2(2,3)(PERCISION) & MULTS_1_9_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_9_3(2,3)(PERCISION) & MULTS_1_9_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(2,3)<=signed(MULTS_1_10_2(2,3)(PERCISION) & MULTS_1_10_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_10_3(2,3)(PERCISION) & MULTS_1_10_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(2,3)<=signed(MULTS_1_11_2(2,3)(PERCISION) & MULTS_1_11_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_11_3(2,3)(PERCISION) & MULTS_1_11_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(2,3)<=signed(MULTS_1_12_2(2,3)(PERCISION) & MULTS_1_12_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_12_3(2,3)(PERCISION) & MULTS_1_12_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(2,3)<=signed(MULTS_1_13_2(2,3)(PERCISION) & MULTS_1_13_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_13_3(2,3)(PERCISION) & MULTS_1_13_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(2,3)<=signed(MULTS_1_14_2(2,3)(PERCISION) & MULTS_1_14_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_14_3(2,3)(PERCISION) & MULTS_1_14_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(2,3)<=signed(MULTS_1_15_2(2,3)(PERCISION) & MULTS_1_15_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_15_3(2,3)(PERCISION) & MULTS_1_15_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(2,3)<=signed(MULTS_1_16_2(2,3)(PERCISION) & MULTS_1_16_2(2,3)(PERCISION downto 1)) + signed(MULTS_1_16_3(2,3)(PERCISION) & MULTS_1_16_3(2,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(2,3) ------------------

			MULTS_2_1_2(2,4)<=signed(MULTS_1_1_2(2,4)(PERCISION) & MULTS_1_1_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_1_3(2,4)(PERCISION) & MULTS_1_1_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(2,4)<=signed(MULTS_1_2_2(2,4)(PERCISION) & MULTS_1_2_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_2_3(2,4)(PERCISION) & MULTS_1_2_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(2,4)<=signed(MULTS_1_3_2(2,4)(PERCISION) & MULTS_1_3_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_3_3(2,4)(PERCISION) & MULTS_1_3_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(2,4)<=signed(MULTS_1_4_2(2,4)(PERCISION) & MULTS_1_4_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_4_3(2,4)(PERCISION) & MULTS_1_4_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(2,4)<=signed(MULTS_1_5_2(2,4)(PERCISION) & MULTS_1_5_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_5_3(2,4)(PERCISION) & MULTS_1_5_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(2,4)<=signed(MULTS_1_6_2(2,4)(PERCISION) & MULTS_1_6_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_6_3(2,4)(PERCISION) & MULTS_1_6_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(2,4)<=signed(MULTS_1_7_2(2,4)(PERCISION) & MULTS_1_7_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_7_3(2,4)(PERCISION) & MULTS_1_7_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(2,4)<=signed(MULTS_1_8_2(2,4)(PERCISION) & MULTS_1_8_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_8_3(2,4)(PERCISION) & MULTS_1_8_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(2,4)<=signed(MULTS_1_9_2(2,4)(PERCISION) & MULTS_1_9_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_9_3(2,4)(PERCISION) & MULTS_1_9_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(2,4)<=signed(MULTS_1_10_2(2,4)(PERCISION) & MULTS_1_10_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_10_3(2,4)(PERCISION) & MULTS_1_10_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(2,4)<=signed(MULTS_1_11_2(2,4)(PERCISION) & MULTS_1_11_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_11_3(2,4)(PERCISION) & MULTS_1_11_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(2,4)<=signed(MULTS_1_12_2(2,4)(PERCISION) & MULTS_1_12_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_12_3(2,4)(PERCISION) & MULTS_1_12_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(2,4)<=signed(MULTS_1_13_2(2,4)(PERCISION) & MULTS_1_13_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_13_3(2,4)(PERCISION) & MULTS_1_13_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(2,4)<=signed(MULTS_1_14_2(2,4)(PERCISION) & MULTS_1_14_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_14_3(2,4)(PERCISION) & MULTS_1_14_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(2,4)<=signed(MULTS_1_15_2(2,4)(PERCISION) & MULTS_1_15_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_15_3(2,4)(PERCISION) & MULTS_1_15_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(2,4)<=signed(MULTS_1_16_2(2,4)(PERCISION) & MULTS_1_16_2(2,4)(PERCISION downto 1)) + signed(MULTS_1_16_3(2,4)(PERCISION) & MULTS_1_16_3(2,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(2,4) ------------------

			MULTS_2_1_2(3,0)<=signed(MULTS_1_1_2(3,0)(PERCISION) & MULTS_1_1_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_1_3(3,0)(PERCISION) & MULTS_1_1_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(3,0)<=signed(MULTS_1_2_2(3,0)(PERCISION) & MULTS_1_2_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_2_3(3,0)(PERCISION) & MULTS_1_2_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(3,0)<=signed(MULTS_1_3_2(3,0)(PERCISION) & MULTS_1_3_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_3_3(3,0)(PERCISION) & MULTS_1_3_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(3,0)<=signed(MULTS_1_4_2(3,0)(PERCISION) & MULTS_1_4_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_4_3(3,0)(PERCISION) & MULTS_1_4_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(3,0)<=signed(MULTS_1_5_2(3,0)(PERCISION) & MULTS_1_5_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_5_3(3,0)(PERCISION) & MULTS_1_5_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(3,0)<=signed(MULTS_1_6_2(3,0)(PERCISION) & MULTS_1_6_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_6_3(3,0)(PERCISION) & MULTS_1_6_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(3,0)<=signed(MULTS_1_7_2(3,0)(PERCISION) & MULTS_1_7_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_7_3(3,0)(PERCISION) & MULTS_1_7_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(3,0)<=signed(MULTS_1_8_2(3,0)(PERCISION) & MULTS_1_8_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_8_3(3,0)(PERCISION) & MULTS_1_8_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(3,0)<=signed(MULTS_1_9_2(3,0)(PERCISION) & MULTS_1_9_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_9_3(3,0)(PERCISION) & MULTS_1_9_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(3,0)<=signed(MULTS_1_10_2(3,0)(PERCISION) & MULTS_1_10_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_10_3(3,0)(PERCISION) & MULTS_1_10_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(3,0)<=signed(MULTS_1_11_2(3,0)(PERCISION) & MULTS_1_11_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_11_3(3,0)(PERCISION) & MULTS_1_11_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(3,0)<=signed(MULTS_1_12_2(3,0)(PERCISION) & MULTS_1_12_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_12_3(3,0)(PERCISION) & MULTS_1_12_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(3,0)<=signed(MULTS_1_13_2(3,0)(PERCISION) & MULTS_1_13_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_13_3(3,0)(PERCISION) & MULTS_1_13_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(3,0)<=signed(MULTS_1_14_2(3,0)(PERCISION) & MULTS_1_14_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_14_3(3,0)(PERCISION) & MULTS_1_14_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(3,0)<=signed(MULTS_1_15_2(3,0)(PERCISION) & MULTS_1_15_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_15_3(3,0)(PERCISION) & MULTS_1_15_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(3,0)<=signed(MULTS_1_16_2(3,0)(PERCISION) & MULTS_1_16_2(3,0)(PERCISION downto 1)) + signed(MULTS_1_16_3(3,0)(PERCISION) & MULTS_1_16_3(3,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(3,0) ------------------

			MULTS_2_1_2(3,1)<=signed(MULTS_1_1_2(3,1)(PERCISION) & MULTS_1_1_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_1_3(3,1)(PERCISION) & MULTS_1_1_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(3,1)<=signed(MULTS_1_2_2(3,1)(PERCISION) & MULTS_1_2_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_2_3(3,1)(PERCISION) & MULTS_1_2_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(3,1)<=signed(MULTS_1_3_2(3,1)(PERCISION) & MULTS_1_3_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_3_3(3,1)(PERCISION) & MULTS_1_3_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(3,1)<=signed(MULTS_1_4_2(3,1)(PERCISION) & MULTS_1_4_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_4_3(3,1)(PERCISION) & MULTS_1_4_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(3,1)<=signed(MULTS_1_5_2(3,1)(PERCISION) & MULTS_1_5_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_5_3(3,1)(PERCISION) & MULTS_1_5_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(3,1)<=signed(MULTS_1_6_2(3,1)(PERCISION) & MULTS_1_6_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_6_3(3,1)(PERCISION) & MULTS_1_6_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(3,1)<=signed(MULTS_1_7_2(3,1)(PERCISION) & MULTS_1_7_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_7_3(3,1)(PERCISION) & MULTS_1_7_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(3,1)<=signed(MULTS_1_8_2(3,1)(PERCISION) & MULTS_1_8_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_8_3(3,1)(PERCISION) & MULTS_1_8_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(3,1)<=signed(MULTS_1_9_2(3,1)(PERCISION) & MULTS_1_9_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_9_3(3,1)(PERCISION) & MULTS_1_9_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(3,1)<=signed(MULTS_1_10_2(3,1)(PERCISION) & MULTS_1_10_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_10_3(3,1)(PERCISION) & MULTS_1_10_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(3,1)<=signed(MULTS_1_11_2(3,1)(PERCISION) & MULTS_1_11_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_11_3(3,1)(PERCISION) & MULTS_1_11_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(3,1)<=signed(MULTS_1_12_2(3,1)(PERCISION) & MULTS_1_12_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_12_3(3,1)(PERCISION) & MULTS_1_12_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(3,1)<=signed(MULTS_1_13_2(3,1)(PERCISION) & MULTS_1_13_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_13_3(3,1)(PERCISION) & MULTS_1_13_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(3,1)<=signed(MULTS_1_14_2(3,1)(PERCISION) & MULTS_1_14_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_14_3(3,1)(PERCISION) & MULTS_1_14_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(3,1)<=signed(MULTS_1_15_2(3,1)(PERCISION) & MULTS_1_15_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_15_3(3,1)(PERCISION) & MULTS_1_15_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(3,1)<=signed(MULTS_1_16_2(3,1)(PERCISION) & MULTS_1_16_2(3,1)(PERCISION downto 1)) + signed(MULTS_1_16_3(3,1)(PERCISION) & MULTS_1_16_3(3,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(3,1) ------------------

			MULTS_2_1_2(3,2)<=signed(MULTS_1_1_2(3,2)(PERCISION) & MULTS_1_1_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_1_3(3,2)(PERCISION) & MULTS_1_1_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(3,2)<=signed(MULTS_1_2_2(3,2)(PERCISION) & MULTS_1_2_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_2_3(3,2)(PERCISION) & MULTS_1_2_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(3,2)<=signed(MULTS_1_3_2(3,2)(PERCISION) & MULTS_1_3_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_3_3(3,2)(PERCISION) & MULTS_1_3_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(3,2)<=signed(MULTS_1_4_2(3,2)(PERCISION) & MULTS_1_4_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_4_3(3,2)(PERCISION) & MULTS_1_4_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(3,2)<=signed(MULTS_1_5_2(3,2)(PERCISION) & MULTS_1_5_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_5_3(3,2)(PERCISION) & MULTS_1_5_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(3,2)<=signed(MULTS_1_6_2(3,2)(PERCISION) & MULTS_1_6_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_6_3(3,2)(PERCISION) & MULTS_1_6_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(3,2)<=signed(MULTS_1_7_2(3,2)(PERCISION) & MULTS_1_7_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_7_3(3,2)(PERCISION) & MULTS_1_7_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(3,2)<=signed(MULTS_1_8_2(3,2)(PERCISION) & MULTS_1_8_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_8_3(3,2)(PERCISION) & MULTS_1_8_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(3,2)<=signed(MULTS_1_9_2(3,2)(PERCISION) & MULTS_1_9_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_9_3(3,2)(PERCISION) & MULTS_1_9_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(3,2)<=signed(MULTS_1_10_2(3,2)(PERCISION) & MULTS_1_10_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_10_3(3,2)(PERCISION) & MULTS_1_10_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(3,2)<=signed(MULTS_1_11_2(3,2)(PERCISION) & MULTS_1_11_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_11_3(3,2)(PERCISION) & MULTS_1_11_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(3,2)<=signed(MULTS_1_12_2(3,2)(PERCISION) & MULTS_1_12_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_12_3(3,2)(PERCISION) & MULTS_1_12_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(3,2)<=signed(MULTS_1_13_2(3,2)(PERCISION) & MULTS_1_13_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_13_3(3,2)(PERCISION) & MULTS_1_13_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(3,2)<=signed(MULTS_1_14_2(3,2)(PERCISION) & MULTS_1_14_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_14_3(3,2)(PERCISION) & MULTS_1_14_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(3,2)<=signed(MULTS_1_15_2(3,2)(PERCISION) & MULTS_1_15_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_15_3(3,2)(PERCISION) & MULTS_1_15_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(3,2)<=signed(MULTS_1_16_2(3,2)(PERCISION) & MULTS_1_16_2(3,2)(PERCISION downto 1)) + signed(MULTS_1_16_3(3,2)(PERCISION) & MULTS_1_16_3(3,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(3,2) ------------------

			MULTS_2_1_2(3,3)<=signed(MULTS_1_1_2(3,3)(PERCISION) & MULTS_1_1_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_1_3(3,3)(PERCISION) & MULTS_1_1_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(3,3)<=signed(MULTS_1_2_2(3,3)(PERCISION) & MULTS_1_2_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_2_3(3,3)(PERCISION) & MULTS_1_2_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(3,3)<=signed(MULTS_1_3_2(3,3)(PERCISION) & MULTS_1_3_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_3_3(3,3)(PERCISION) & MULTS_1_3_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(3,3)<=signed(MULTS_1_4_2(3,3)(PERCISION) & MULTS_1_4_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_4_3(3,3)(PERCISION) & MULTS_1_4_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(3,3)<=signed(MULTS_1_5_2(3,3)(PERCISION) & MULTS_1_5_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_5_3(3,3)(PERCISION) & MULTS_1_5_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(3,3)<=signed(MULTS_1_6_2(3,3)(PERCISION) & MULTS_1_6_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_6_3(3,3)(PERCISION) & MULTS_1_6_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(3,3)<=signed(MULTS_1_7_2(3,3)(PERCISION) & MULTS_1_7_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_7_3(3,3)(PERCISION) & MULTS_1_7_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(3,3)<=signed(MULTS_1_8_2(3,3)(PERCISION) & MULTS_1_8_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_8_3(3,3)(PERCISION) & MULTS_1_8_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(3,3)<=signed(MULTS_1_9_2(3,3)(PERCISION) & MULTS_1_9_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_9_3(3,3)(PERCISION) & MULTS_1_9_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(3,3)<=signed(MULTS_1_10_2(3,3)(PERCISION) & MULTS_1_10_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_10_3(3,3)(PERCISION) & MULTS_1_10_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(3,3)<=signed(MULTS_1_11_2(3,3)(PERCISION) & MULTS_1_11_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_11_3(3,3)(PERCISION) & MULTS_1_11_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(3,3)<=signed(MULTS_1_12_2(3,3)(PERCISION) & MULTS_1_12_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_12_3(3,3)(PERCISION) & MULTS_1_12_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(3,3)<=signed(MULTS_1_13_2(3,3)(PERCISION) & MULTS_1_13_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_13_3(3,3)(PERCISION) & MULTS_1_13_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(3,3)<=signed(MULTS_1_14_2(3,3)(PERCISION) & MULTS_1_14_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_14_3(3,3)(PERCISION) & MULTS_1_14_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(3,3)<=signed(MULTS_1_15_2(3,3)(PERCISION) & MULTS_1_15_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_15_3(3,3)(PERCISION) & MULTS_1_15_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(3,3)<=signed(MULTS_1_16_2(3,3)(PERCISION) & MULTS_1_16_2(3,3)(PERCISION downto 1)) + signed(MULTS_1_16_3(3,3)(PERCISION) & MULTS_1_16_3(3,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(3,3) ------------------

			MULTS_2_1_2(3,4)<=signed(MULTS_1_1_2(3,4)(PERCISION) & MULTS_1_1_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_1_3(3,4)(PERCISION) & MULTS_1_1_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(3,4)<=signed(MULTS_1_2_2(3,4)(PERCISION) & MULTS_1_2_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_2_3(3,4)(PERCISION) & MULTS_1_2_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(3,4)<=signed(MULTS_1_3_2(3,4)(PERCISION) & MULTS_1_3_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_3_3(3,4)(PERCISION) & MULTS_1_3_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(3,4)<=signed(MULTS_1_4_2(3,4)(PERCISION) & MULTS_1_4_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_4_3(3,4)(PERCISION) & MULTS_1_4_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(3,4)<=signed(MULTS_1_5_2(3,4)(PERCISION) & MULTS_1_5_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_5_3(3,4)(PERCISION) & MULTS_1_5_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(3,4)<=signed(MULTS_1_6_2(3,4)(PERCISION) & MULTS_1_6_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_6_3(3,4)(PERCISION) & MULTS_1_6_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(3,4)<=signed(MULTS_1_7_2(3,4)(PERCISION) & MULTS_1_7_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_7_3(3,4)(PERCISION) & MULTS_1_7_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(3,4)<=signed(MULTS_1_8_2(3,4)(PERCISION) & MULTS_1_8_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_8_3(3,4)(PERCISION) & MULTS_1_8_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(3,4)<=signed(MULTS_1_9_2(3,4)(PERCISION) & MULTS_1_9_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_9_3(3,4)(PERCISION) & MULTS_1_9_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(3,4)<=signed(MULTS_1_10_2(3,4)(PERCISION) & MULTS_1_10_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_10_3(3,4)(PERCISION) & MULTS_1_10_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(3,4)<=signed(MULTS_1_11_2(3,4)(PERCISION) & MULTS_1_11_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_11_3(3,4)(PERCISION) & MULTS_1_11_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(3,4)<=signed(MULTS_1_12_2(3,4)(PERCISION) & MULTS_1_12_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_12_3(3,4)(PERCISION) & MULTS_1_12_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(3,4)<=signed(MULTS_1_13_2(3,4)(PERCISION) & MULTS_1_13_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_13_3(3,4)(PERCISION) & MULTS_1_13_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(3,4)<=signed(MULTS_1_14_2(3,4)(PERCISION) & MULTS_1_14_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_14_3(3,4)(PERCISION) & MULTS_1_14_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(3,4)<=signed(MULTS_1_15_2(3,4)(PERCISION) & MULTS_1_15_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_15_3(3,4)(PERCISION) & MULTS_1_15_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(3,4)<=signed(MULTS_1_16_2(3,4)(PERCISION) & MULTS_1_16_2(3,4)(PERCISION downto 1)) + signed(MULTS_1_16_3(3,4)(PERCISION) & MULTS_1_16_3(3,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(3,4) ------------------

			MULTS_2_1_2(4,0)<=signed(MULTS_1_1_2(4,0)(PERCISION) & MULTS_1_1_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_1_3(4,0)(PERCISION) & MULTS_1_1_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(4,0)<=signed(MULTS_1_2_2(4,0)(PERCISION) & MULTS_1_2_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_2_3(4,0)(PERCISION) & MULTS_1_2_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(4,0)<=signed(MULTS_1_3_2(4,0)(PERCISION) & MULTS_1_3_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_3_3(4,0)(PERCISION) & MULTS_1_3_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(4,0)<=signed(MULTS_1_4_2(4,0)(PERCISION) & MULTS_1_4_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_4_3(4,0)(PERCISION) & MULTS_1_4_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(4,0)<=signed(MULTS_1_5_2(4,0)(PERCISION) & MULTS_1_5_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_5_3(4,0)(PERCISION) & MULTS_1_5_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(4,0)<=signed(MULTS_1_6_2(4,0)(PERCISION) & MULTS_1_6_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_6_3(4,0)(PERCISION) & MULTS_1_6_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(4,0)<=signed(MULTS_1_7_2(4,0)(PERCISION) & MULTS_1_7_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_7_3(4,0)(PERCISION) & MULTS_1_7_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(4,0)<=signed(MULTS_1_8_2(4,0)(PERCISION) & MULTS_1_8_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_8_3(4,0)(PERCISION) & MULTS_1_8_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(4,0)<=signed(MULTS_1_9_2(4,0)(PERCISION) & MULTS_1_9_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_9_3(4,0)(PERCISION) & MULTS_1_9_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(4,0)<=signed(MULTS_1_10_2(4,0)(PERCISION) & MULTS_1_10_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_10_3(4,0)(PERCISION) & MULTS_1_10_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(4,0)<=signed(MULTS_1_11_2(4,0)(PERCISION) & MULTS_1_11_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_11_3(4,0)(PERCISION) & MULTS_1_11_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(4,0)<=signed(MULTS_1_12_2(4,0)(PERCISION) & MULTS_1_12_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_12_3(4,0)(PERCISION) & MULTS_1_12_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(4,0)<=signed(MULTS_1_13_2(4,0)(PERCISION) & MULTS_1_13_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_13_3(4,0)(PERCISION) & MULTS_1_13_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(4,0)<=signed(MULTS_1_14_2(4,0)(PERCISION) & MULTS_1_14_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_14_3(4,0)(PERCISION) & MULTS_1_14_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(4,0)<=signed(MULTS_1_15_2(4,0)(PERCISION) & MULTS_1_15_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_15_3(4,0)(PERCISION) & MULTS_1_15_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(4,0)<=signed(MULTS_1_16_2(4,0)(PERCISION) & MULTS_1_16_2(4,0)(PERCISION downto 1)) + signed(MULTS_1_16_3(4,0)(PERCISION) & MULTS_1_16_3(4,0)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(4,0) ------------------

			MULTS_2_1_2(4,1)<=signed(MULTS_1_1_2(4,1)(PERCISION) & MULTS_1_1_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_1_3(4,1)(PERCISION) & MULTS_1_1_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(4,1)<=signed(MULTS_1_2_2(4,1)(PERCISION) & MULTS_1_2_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_2_3(4,1)(PERCISION) & MULTS_1_2_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(4,1)<=signed(MULTS_1_3_2(4,1)(PERCISION) & MULTS_1_3_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_3_3(4,1)(PERCISION) & MULTS_1_3_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(4,1)<=signed(MULTS_1_4_2(4,1)(PERCISION) & MULTS_1_4_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_4_3(4,1)(PERCISION) & MULTS_1_4_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(4,1)<=signed(MULTS_1_5_2(4,1)(PERCISION) & MULTS_1_5_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_5_3(4,1)(PERCISION) & MULTS_1_5_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(4,1)<=signed(MULTS_1_6_2(4,1)(PERCISION) & MULTS_1_6_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_6_3(4,1)(PERCISION) & MULTS_1_6_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(4,1)<=signed(MULTS_1_7_2(4,1)(PERCISION) & MULTS_1_7_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_7_3(4,1)(PERCISION) & MULTS_1_7_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(4,1)<=signed(MULTS_1_8_2(4,1)(PERCISION) & MULTS_1_8_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_8_3(4,1)(PERCISION) & MULTS_1_8_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(4,1)<=signed(MULTS_1_9_2(4,1)(PERCISION) & MULTS_1_9_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_9_3(4,1)(PERCISION) & MULTS_1_9_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(4,1)<=signed(MULTS_1_10_2(4,1)(PERCISION) & MULTS_1_10_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_10_3(4,1)(PERCISION) & MULTS_1_10_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(4,1)<=signed(MULTS_1_11_2(4,1)(PERCISION) & MULTS_1_11_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_11_3(4,1)(PERCISION) & MULTS_1_11_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(4,1)<=signed(MULTS_1_12_2(4,1)(PERCISION) & MULTS_1_12_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_12_3(4,1)(PERCISION) & MULTS_1_12_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(4,1)<=signed(MULTS_1_13_2(4,1)(PERCISION) & MULTS_1_13_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_13_3(4,1)(PERCISION) & MULTS_1_13_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(4,1)<=signed(MULTS_1_14_2(4,1)(PERCISION) & MULTS_1_14_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_14_3(4,1)(PERCISION) & MULTS_1_14_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(4,1)<=signed(MULTS_1_15_2(4,1)(PERCISION) & MULTS_1_15_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_15_3(4,1)(PERCISION) & MULTS_1_15_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(4,1)<=signed(MULTS_1_16_2(4,1)(PERCISION) & MULTS_1_16_2(4,1)(PERCISION downto 1)) + signed(MULTS_1_16_3(4,1)(PERCISION) & MULTS_1_16_3(4,1)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(4,1) ------------------

			MULTS_2_1_2(4,2)<=signed(MULTS_1_1_2(4,2)(PERCISION) & MULTS_1_1_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_1_3(4,2)(PERCISION) & MULTS_1_1_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(4,2)<=signed(MULTS_1_2_2(4,2)(PERCISION) & MULTS_1_2_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_2_3(4,2)(PERCISION) & MULTS_1_2_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(4,2)<=signed(MULTS_1_3_2(4,2)(PERCISION) & MULTS_1_3_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_3_3(4,2)(PERCISION) & MULTS_1_3_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(4,2)<=signed(MULTS_1_4_2(4,2)(PERCISION) & MULTS_1_4_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_4_3(4,2)(PERCISION) & MULTS_1_4_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(4,2)<=signed(MULTS_1_5_2(4,2)(PERCISION) & MULTS_1_5_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_5_3(4,2)(PERCISION) & MULTS_1_5_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(4,2)<=signed(MULTS_1_6_2(4,2)(PERCISION) & MULTS_1_6_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_6_3(4,2)(PERCISION) & MULTS_1_6_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(4,2)<=signed(MULTS_1_7_2(4,2)(PERCISION) & MULTS_1_7_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_7_3(4,2)(PERCISION) & MULTS_1_7_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(4,2)<=signed(MULTS_1_8_2(4,2)(PERCISION) & MULTS_1_8_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_8_3(4,2)(PERCISION) & MULTS_1_8_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(4,2)<=signed(MULTS_1_9_2(4,2)(PERCISION) & MULTS_1_9_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_9_3(4,2)(PERCISION) & MULTS_1_9_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(4,2)<=signed(MULTS_1_10_2(4,2)(PERCISION) & MULTS_1_10_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_10_3(4,2)(PERCISION) & MULTS_1_10_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(4,2)<=signed(MULTS_1_11_2(4,2)(PERCISION) & MULTS_1_11_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_11_3(4,2)(PERCISION) & MULTS_1_11_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(4,2)<=signed(MULTS_1_12_2(4,2)(PERCISION) & MULTS_1_12_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_12_3(4,2)(PERCISION) & MULTS_1_12_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(4,2)<=signed(MULTS_1_13_2(4,2)(PERCISION) & MULTS_1_13_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_13_3(4,2)(PERCISION) & MULTS_1_13_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(4,2)<=signed(MULTS_1_14_2(4,2)(PERCISION) & MULTS_1_14_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_14_3(4,2)(PERCISION) & MULTS_1_14_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(4,2)<=signed(MULTS_1_15_2(4,2)(PERCISION) & MULTS_1_15_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_15_3(4,2)(PERCISION) & MULTS_1_15_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(4,2)<=signed(MULTS_1_16_2(4,2)(PERCISION) & MULTS_1_16_2(4,2)(PERCISION downto 1)) + signed(MULTS_1_16_3(4,2)(PERCISION) & MULTS_1_16_3(4,2)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(4,2) ------------------

			MULTS_2_1_2(4,3)<=signed(MULTS_1_1_2(4,3)(PERCISION) & MULTS_1_1_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_1_3(4,3)(PERCISION) & MULTS_1_1_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(4,3)<=signed(MULTS_1_2_2(4,3)(PERCISION) & MULTS_1_2_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_2_3(4,3)(PERCISION) & MULTS_1_2_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(4,3)<=signed(MULTS_1_3_2(4,3)(PERCISION) & MULTS_1_3_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_3_3(4,3)(PERCISION) & MULTS_1_3_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(4,3)<=signed(MULTS_1_4_2(4,3)(PERCISION) & MULTS_1_4_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_4_3(4,3)(PERCISION) & MULTS_1_4_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(4,3)<=signed(MULTS_1_5_2(4,3)(PERCISION) & MULTS_1_5_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_5_3(4,3)(PERCISION) & MULTS_1_5_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(4,3)<=signed(MULTS_1_6_2(4,3)(PERCISION) & MULTS_1_6_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_6_3(4,3)(PERCISION) & MULTS_1_6_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(4,3)<=signed(MULTS_1_7_2(4,3)(PERCISION) & MULTS_1_7_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_7_3(4,3)(PERCISION) & MULTS_1_7_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(4,3)<=signed(MULTS_1_8_2(4,3)(PERCISION) & MULTS_1_8_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_8_3(4,3)(PERCISION) & MULTS_1_8_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(4,3)<=signed(MULTS_1_9_2(4,3)(PERCISION) & MULTS_1_9_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_9_3(4,3)(PERCISION) & MULTS_1_9_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(4,3)<=signed(MULTS_1_10_2(4,3)(PERCISION) & MULTS_1_10_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_10_3(4,3)(PERCISION) & MULTS_1_10_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(4,3)<=signed(MULTS_1_11_2(4,3)(PERCISION) & MULTS_1_11_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_11_3(4,3)(PERCISION) & MULTS_1_11_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(4,3)<=signed(MULTS_1_12_2(4,3)(PERCISION) & MULTS_1_12_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_12_3(4,3)(PERCISION) & MULTS_1_12_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(4,3)<=signed(MULTS_1_13_2(4,3)(PERCISION) & MULTS_1_13_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_13_3(4,3)(PERCISION) & MULTS_1_13_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(4,3)<=signed(MULTS_1_14_2(4,3)(PERCISION) & MULTS_1_14_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_14_3(4,3)(PERCISION) & MULTS_1_14_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(4,3)<=signed(MULTS_1_15_2(4,3)(PERCISION) & MULTS_1_15_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_15_3(4,3)(PERCISION) & MULTS_1_15_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(4,3)<=signed(MULTS_1_16_2(4,3)(PERCISION) & MULTS_1_16_2(4,3)(PERCISION downto 1)) + signed(MULTS_1_16_3(4,3)(PERCISION) & MULTS_1_16_3(4,3)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(4,3) ------------------

			MULTS_2_1_2(4,4)<=signed(MULTS_1_1_2(4,4)(PERCISION) & MULTS_1_1_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_1_3(4,4)(PERCISION) & MULTS_1_1_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(1) ------------------

			MULTS_2_2_2(4,4)<=signed(MULTS_1_2_2(4,4)(PERCISION) & MULTS_1_2_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_2_3(4,4)(PERCISION) & MULTS_1_2_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(2) ------------------

			MULTS_2_3_2(4,4)<=signed(MULTS_1_3_2(4,4)(PERCISION) & MULTS_1_3_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_3_3(4,4)(PERCISION) & MULTS_1_3_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(3) ------------------

			MULTS_2_4_2(4,4)<=signed(MULTS_1_4_2(4,4)(PERCISION) & MULTS_1_4_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_4_3(4,4)(PERCISION) & MULTS_1_4_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(4) ------------------

			MULTS_2_5_2(4,4)<=signed(MULTS_1_5_2(4,4)(PERCISION) & MULTS_1_5_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_5_3(4,4)(PERCISION) & MULTS_1_5_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(5) ------------------

			MULTS_2_6_2(4,4)<=signed(MULTS_1_6_2(4,4)(PERCISION) & MULTS_1_6_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_6_3(4,4)(PERCISION) & MULTS_1_6_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(6) ------------------

			MULTS_2_7_2(4,4)<=signed(MULTS_1_7_2(4,4)(PERCISION) & MULTS_1_7_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_7_3(4,4)(PERCISION) & MULTS_1_7_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(7) ------------------

			MULTS_2_8_2(4,4)<=signed(MULTS_1_8_2(4,4)(PERCISION) & MULTS_1_8_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_8_3(4,4)(PERCISION) & MULTS_1_8_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(8) ------------------

			MULTS_2_9_2(4,4)<=signed(MULTS_1_9_2(4,4)(PERCISION) & MULTS_1_9_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_9_3(4,4)(PERCISION) & MULTS_1_9_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(9) ------------------

			MULTS_2_10_2(4,4)<=signed(MULTS_1_10_2(4,4)(PERCISION) & MULTS_1_10_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_10_3(4,4)(PERCISION) & MULTS_1_10_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(10) ------------------

			MULTS_2_11_2(4,4)<=signed(MULTS_1_11_2(4,4)(PERCISION) & MULTS_1_11_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_11_3(4,4)(PERCISION) & MULTS_1_11_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(11) ------------------

			MULTS_2_12_2(4,4)<=signed(MULTS_1_12_2(4,4)(PERCISION) & MULTS_1_12_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_12_3(4,4)(PERCISION) & MULTS_1_12_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(12) ------------------

			MULTS_2_13_2(4,4)<=signed(MULTS_1_13_2(4,4)(PERCISION) & MULTS_1_13_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_13_3(4,4)(PERCISION) & MULTS_1_13_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(13) ------------------

			MULTS_2_14_2(4,4)<=signed(MULTS_1_14_2(4,4)(PERCISION) & MULTS_1_14_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_14_3(4,4)(PERCISION) & MULTS_1_14_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(14) ------------------

			MULTS_2_15_2(4,4)<=signed(MULTS_1_15_2(4,4)(PERCISION) & MULTS_1_15_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_15_3(4,4)(PERCISION) & MULTS_1_15_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(15) ------------------

			MULTS_2_16_2(4,4)<=signed(MULTS_1_16_2(4,4)(PERCISION) & MULTS_1_16_2(4,4)(PERCISION downto 1)) + signed(MULTS_1_16_3(4,4)(PERCISION) & MULTS_1_16_3(4,4)(PERCISION downto 1));
                        ---------------------SUM P_MAPS of FMAP(16) ------------------

                            -----------------------END OF INDEX(4,4) ------------------



                     EN_SUM_MULT_3<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_3 = '1' then
			------------------------------------STAGE-3--------------------------------------
			MULTS_3_1_1(0,0)<=signed(MULTS_2_1_1(0,0)(PERCISION) & MULTS_2_1_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_1_2(0,0)(PERCISION) & MULTS_2_1_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(0,0)<=signed(MULTS_2_2_1(0,0)(PERCISION) & MULTS_2_2_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_2_2(0,0)(PERCISION) & MULTS_2_2_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(0,0)<=signed(MULTS_2_3_1(0,0)(PERCISION) & MULTS_2_3_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_3_2(0,0)(PERCISION) & MULTS_2_3_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(0,0)<=signed(MULTS_2_4_1(0,0)(PERCISION) & MULTS_2_4_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_4_2(0,0)(PERCISION) & MULTS_2_4_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(0,0)<=signed(MULTS_2_5_1(0,0)(PERCISION) & MULTS_2_5_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_5_2(0,0)(PERCISION) & MULTS_2_5_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(0,0)<=signed(MULTS_2_6_1(0,0)(PERCISION) & MULTS_2_6_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_6_2(0,0)(PERCISION) & MULTS_2_6_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(0,0)<=signed(MULTS_2_7_1(0,0)(PERCISION) & MULTS_2_7_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_7_2(0,0)(PERCISION) & MULTS_2_7_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(0,0)<=signed(MULTS_2_8_1(0,0)(PERCISION) & MULTS_2_8_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_8_2(0,0)(PERCISION) & MULTS_2_8_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(0,0)<=signed(MULTS_2_9_1(0,0)(PERCISION) & MULTS_2_9_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_9_2(0,0)(PERCISION) & MULTS_2_9_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(0,0)<=signed(MULTS_2_10_1(0,0)(PERCISION) & MULTS_2_10_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_10_2(0,0)(PERCISION) & MULTS_2_10_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(0,0)<=signed(MULTS_2_11_1(0,0)(PERCISION) & MULTS_2_11_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_11_2(0,0)(PERCISION) & MULTS_2_11_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(0,0)<=signed(MULTS_2_12_1(0,0)(PERCISION) & MULTS_2_12_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_12_2(0,0)(PERCISION) & MULTS_2_12_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(0,0)<=signed(MULTS_2_13_1(0,0)(PERCISION) & MULTS_2_13_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_13_2(0,0)(PERCISION) & MULTS_2_13_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(0,0)<=signed(MULTS_2_14_1(0,0)(PERCISION) & MULTS_2_14_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_14_2(0,0)(PERCISION) & MULTS_2_14_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(0,0)<=signed(MULTS_2_15_1(0,0)(PERCISION) & MULTS_2_15_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_15_2(0,0)(PERCISION) & MULTS_2_15_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(0,0)<=signed(MULTS_2_16_1(0,0)(PERCISION) & MULTS_2_16_1(0,0)(PERCISION downto 1)) + signed(MULTS_2_16_2(0,0)(PERCISION) & MULTS_2_16_2(0,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(0,0) ------------------

			MULTS_3_1_1(0,1)<=signed(MULTS_2_1_1(0,1)(PERCISION) & MULTS_2_1_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_1_2(0,1)(PERCISION) & MULTS_2_1_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(0,1)<=signed(MULTS_2_2_1(0,1)(PERCISION) & MULTS_2_2_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_2_2(0,1)(PERCISION) & MULTS_2_2_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(0,1)<=signed(MULTS_2_3_1(0,1)(PERCISION) & MULTS_2_3_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_3_2(0,1)(PERCISION) & MULTS_2_3_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(0,1)<=signed(MULTS_2_4_1(0,1)(PERCISION) & MULTS_2_4_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_4_2(0,1)(PERCISION) & MULTS_2_4_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(0,1)<=signed(MULTS_2_5_1(0,1)(PERCISION) & MULTS_2_5_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_5_2(0,1)(PERCISION) & MULTS_2_5_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(0,1)<=signed(MULTS_2_6_1(0,1)(PERCISION) & MULTS_2_6_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_6_2(0,1)(PERCISION) & MULTS_2_6_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(0,1)<=signed(MULTS_2_7_1(0,1)(PERCISION) & MULTS_2_7_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_7_2(0,1)(PERCISION) & MULTS_2_7_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(0,1)<=signed(MULTS_2_8_1(0,1)(PERCISION) & MULTS_2_8_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_8_2(0,1)(PERCISION) & MULTS_2_8_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(0,1)<=signed(MULTS_2_9_1(0,1)(PERCISION) & MULTS_2_9_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_9_2(0,1)(PERCISION) & MULTS_2_9_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(0,1)<=signed(MULTS_2_10_1(0,1)(PERCISION) & MULTS_2_10_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_10_2(0,1)(PERCISION) & MULTS_2_10_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(0,1)<=signed(MULTS_2_11_1(0,1)(PERCISION) & MULTS_2_11_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_11_2(0,1)(PERCISION) & MULTS_2_11_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(0,1)<=signed(MULTS_2_12_1(0,1)(PERCISION) & MULTS_2_12_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_12_2(0,1)(PERCISION) & MULTS_2_12_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(0,1)<=signed(MULTS_2_13_1(0,1)(PERCISION) & MULTS_2_13_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_13_2(0,1)(PERCISION) & MULTS_2_13_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(0,1)<=signed(MULTS_2_14_1(0,1)(PERCISION) & MULTS_2_14_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_14_2(0,1)(PERCISION) & MULTS_2_14_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(0,1)<=signed(MULTS_2_15_1(0,1)(PERCISION) & MULTS_2_15_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_15_2(0,1)(PERCISION) & MULTS_2_15_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(0,1)<=signed(MULTS_2_16_1(0,1)(PERCISION) & MULTS_2_16_1(0,1)(PERCISION downto 1)) + signed(MULTS_2_16_2(0,1)(PERCISION) & MULTS_2_16_2(0,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(0,1) ------------------

			MULTS_3_1_1(0,2)<=signed(MULTS_2_1_1(0,2)(PERCISION) & MULTS_2_1_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_1_2(0,2)(PERCISION) & MULTS_2_1_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(0,2)<=signed(MULTS_2_2_1(0,2)(PERCISION) & MULTS_2_2_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_2_2(0,2)(PERCISION) & MULTS_2_2_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(0,2)<=signed(MULTS_2_3_1(0,2)(PERCISION) & MULTS_2_3_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_3_2(0,2)(PERCISION) & MULTS_2_3_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(0,2)<=signed(MULTS_2_4_1(0,2)(PERCISION) & MULTS_2_4_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_4_2(0,2)(PERCISION) & MULTS_2_4_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(0,2)<=signed(MULTS_2_5_1(0,2)(PERCISION) & MULTS_2_5_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_5_2(0,2)(PERCISION) & MULTS_2_5_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(0,2)<=signed(MULTS_2_6_1(0,2)(PERCISION) & MULTS_2_6_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_6_2(0,2)(PERCISION) & MULTS_2_6_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(0,2)<=signed(MULTS_2_7_1(0,2)(PERCISION) & MULTS_2_7_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_7_2(0,2)(PERCISION) & MULTS_2_7_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(0,2)<=signed(MULTS_2_8_1(0,2)(PERCISION) & MULTS_2_8_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_8_2(0,2)(PERCISION) & MULTS_2_8_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(0,2)<=signed(MULTS_2_9_1(0,2)(PERCISION) & MULTS_2_9_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_9_2(0,2)(PERCISION) & MULTS_2_9_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(0,2)<=signed(MULTS_2_10_1(0,2)(PERCISION) & MULTS_2_10_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_10_2(0,2)(PERCISION) & MULTS_2_10_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(0,2)<=signed(MULTS_2_11_1(0,2)(PERCISION) & MULTS_2_11_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_11_2(0,2)(PERCISION) & MULTS_2_11_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(0,2)<=signed(MULTS_2_12_1(0,2)(PERCISION) & MULTS_2_12_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_12_2(0,2)(PERCISION) & MULTS_2_12_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(0,2)<=signed(MULTS_2_13_1(0,2)(PERCISION) & MULTS_2_13_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_13_2(0,2)(PERCISION) & MULTS_2_13_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(0,2)<=signed(MULTS_2_14_1(0,2)(PERCISION) & MULTS_2_14_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_14_2(0,2)(PERCISION) & MULTS_2_14_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(0,2)<=signed(MULTS_2_15_1(0,2)(PERCISION) & MULTS_2_15_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_15_2(0,2)(PERCISION) & MULTS_2_15_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(0,2)<=signed(MULTS_2_16_1(0,2)(PERCISION) & MULTS_2_16_1(0,2)(PERCISION downto 1)) + signed(MULTS_2_16_2(0,2)(PERCISION) & MULTS_2_16_2(0,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(0,2) ------------------

			MULTS_3_1_1(0,3)<=signed(MULTS_2_1_1(0,3)(PERCISION) & MULTS_2_1_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_1_2(0,3)(PERCISION) & MULTS_2_1_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(0,3)<=signed(MULTS_2_2_1(0,3)(PERCISION) & MULTS_2_2_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_2_2(0,3)(PERCISION) & MULTS_2_2_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(0,3)<=signed(MULTS_2_3_1(0,3)(PERCISION) & MULTS_2_3_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_3_2(0,3)(PERCISION) & MULTS_2_3_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(0,3)<=signed(MULTS_2_4_1(0,3)(PERCISION) & MULTS_2_4_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_4_2(0,3)(PERCISION) & MULTS_2_4_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(0,3)<=signed(MULTS_2_5_1(0,3)(PERCISION) & MULTS_2_5_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_5_2(0,3)(PERCISION) & MULTS_2_5_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(0,3)<=signed(MULTS_2_6_1(0,3)(PERCISION) & MULTS_2_6_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_6_2(0,3)(PERCISION) & MULTS_2_6_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(0,3)<=signed(MULTS_2_7_1(0,3)(PERCISION) & MULTS_2_7_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_7_2(0,3)(PERCISION) & MULTS_2_7_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(0,3)<=signed(MULTS_2_8_1(0,3)(PERCISION) & MULTS_2_8_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_8_2(0,3)(PERCISION) & MULTS_2_8_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(0,3)<=signed(MULTS_2_9_1(0,3)(PERCISION) & MULTS_2_9_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_9_2(0,3)(PERCISION) & MULTS_2_9_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(0,3)<=signed(MULTS_2_10_1(0,3)(PERCISION) & MULTS_2_10_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_10_2(0,3)(PERCISION) & MULTS_2_10_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(0,3)<=signed(MULTS_2_11_1(0,3)(PERCISION) & MULTS_2_11_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_11_2(0,3)(PERCISION) & MULTS_2_11_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(0,3)<=signed(MULTS_2_12_1(0,3)(PERCISION) & MULTS_2_12_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_12_2(0,3)(PERCISION) & MULTS_2_12_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(0,3)<=signed(MULTS_2_13_1(0,3)(PERCISION) & MULTS_2_13_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_13_2(0,3)(PERCISION) & MULTS_2_13_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(0,3)<=signed(MULTS_2_14_1(0,3)(PERCISION) & MULTS_2_14_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_14_2(0,3)(PERCISION) & MULTS_2_14_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(0,3)<=signed(MULTS_2_15_1(0,3)(PERCISION) & MULTS_2_15_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_15_2(0,3)(PERCISION) & MULTS_2_15_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(0,3)<=signed(MULTS_2_16_1(0,3)(PERCISION) & MULTS_2_16_1(0,3)(PERCISION downto 1)) + signed(MULTS_2_16_2(0,3)(PERCISION) & MULTS_2_16_2(0,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(0,3) ------------------

			MULTS_3_1_1(0,4)<=signed(MULTS_2_1_1(0,4)(PERCISION) & MULTS_2_1_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_1_2(0,4)(PERCISION) & MULTS_2_1_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(0,4)<=signed(MULTS_2_2_1(0,4)(PERCISION) & MULTS_2_2_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_2_2(0,4)(PERCISION) & MULTS_2_2_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(0,4)<=signed(MULTS_2_3_1(0,4)(PERCISION) & MULTS_2_3_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_3_2(0,4)(PERCISION) & MULTS_2_3_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(0,4)<=signed(MULTS_2_4_1(0,4)(PERCISION) & MULTS_2_4_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_4_2(0,4)(PERCISION) & MULTS_2_4_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(0,4)<=signed(MULTS_2_5_1(0,4)(PERCISION) & MULTS_2_5_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_5_2(0,4)(PERCISION) & MULTS_2_5_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(0,4)<=signed(MULTS_2_6_1(0,4)(PERCISION) & MULTS_2_6_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_6_2(0,4)(PERCISION) & MULTS_2_6_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(0,4)<=signed(MULTS_2_7_1(0,4)(PERCISION) & MULTS_2_7_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_7_2(0,4)(PERCISION) & MULTS_2_7_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(0,4)<=signed(MULTS_2_8_1(0,4)(PERCISION) & MULTS_2_8_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_8_2(0,4)(PERCISION) & MULTS_2_8_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(0,4)<=signed(MULTS_2_9_1(0,4)(PERCISION) & MULTS_2_9_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_9_2(0,4)(PERCISION) & MULTS_2_9_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(0,4)<=signed(MULTS_2_10_1(0,4)(PERCISION) & MULTS_2_10_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_10_2(0,4)(PERCISION) & MULTS_2_10_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(0,4)<=signed(MULTS_2_11_1(0,4)(PERCISION) & MULTS_2_11_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_11_2(0,4)(PERCISION) & MULTS_2_11_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(0,4)<=signed(MULTS_2_12_1(0,4)(PERCISION) & MULTS_2_12_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_12_2(0,4)(PERCISION) & MULTS_2_12_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(0,4)<=signed(MULTS_2_13_1(0,4)(PERCISION) & MULTS_2_13_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_13_2(0,4)(PERCISION) & MULTS_2_13_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(0,4)<=signed(MULTS_2_14_1(0,4)(PERCISION) & MULTS_2_14_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_14_2(0,4)(PERCISION) & MULTS_2_14_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(0,4)<=signed(MULTS_2_15_1(0,4)(PERCISION) & MULTS_2_15_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_15_2(0,4)(PERCISION) & MULTS_2_15_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(0,4)<=signed(MULTS_2_16_1(0,4)(PERCISION) & MULTS_2_16_1(0,4)(PERCISION downto 1)) + signed(MULTS_2_16_2(0,4)(PERCISION) & MULTS_2_16_2(0,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(0,4) ------------------

			MULTS_3_1_1(1,0)<=signed(MULTS_2_1_1(1,0)(PERCISION) & MULTS_2_1_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_1_2(1,0)(PERCISION) & MULTS_2_1_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(1,0)<=signed(MULTS_2_2_1(1,0)(PERCISION) & MULTS_2_2_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_2_2(1,0)(PERCISION) & MULTS_2_2_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(1,0)<=signed(MULTS_2_3_1(1,0)(PERCISION) & MULTS_2_3_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_3_2(1,0)(PERCISION) & MULTS_2_3_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(1,0)<=signed(MULTS_2_4_1(1,0)(PERCISION) & MULTS_2_4_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_4_2(1,0)(PERCISION) & MULTS_2_4_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(1,0)<=signed(MULTS_2_5_1(1,0)(PERCISION) & MULTS_2_5_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_5_2(1,0)(PERCISION) & MULTS_2_5_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(1,0)<=signed(MULTS_2_6_1(1,0)(PERCISION) & MULTS_2_6_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_6_2(1,0)(PERCISION) & MULTS_2_6_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(1,0)<=signed(MULTS_2_7_1(1,0)(PERCISION) & MULTS_2_7_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_7_2(1,0)(PERCISION) & MULTS_2_7_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(1,0)<=signed(MULTS_2_8_1(1,0)(PERCISION) & MULTS_2_8_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_8_2(1,0)(PERCISION) & MULTS_2_8_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(1,0)<=signed(MULTS_2_9_1(1,0)(PERCISION) & MULTS_2_9_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_9_2(1,0)(PERCISION) & MULTS_2_9_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(1,0)<=signed(MULTS_2_10_1(1,0)(PERCISION) & MULTS_2_10_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_10_2(1,0)(PERCISION) & MULTS_2_10_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(1,0)<=signed(MULTS_2_11_1(1,0)(PERCISION) & MULTS_2_11_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_11_2(1,0)(PERCISION) & MULTS_2_11_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(1,0)<=signed(MULTS_2_12_1(1,0)(PERCISION) & MULTS_2_12_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_12_2(1,0)(PERCISION) & MULTS_2_12_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(1,0)<=signed(MULTS_2_13_1(1,0)(PERCISION) & MULTS_2_13_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_13_2(1,0)(PERCISION) & MULTS_2_13_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(1,0)<=signed(MULTS_2_14_1(1,0)(PERCISION) & MULTS_2_14_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_14_2(1,0)(PERCISION) & MULTS_2_14_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(1,0)<=signed(MULTS_2_15_1(1,0)(PERCISION) & MULTS_2_15_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_15_2(1,0)(PERCISION) & MULTS_2_15_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(1,0)<=signed(MULTS_2_16_1(1,0)(PERCISION) & MULTS_2_16_1(1,0)(PERCISION downto 1)) + signed(MULTS_2_16_2(1,0)(PERCISION) & MULTS_2_16_2(1,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(1,0) ------------------

			MULTS_3_1_1(1,1)<=signed(MULTS_2_1_1(1,1)(PERCISION) & MULTS_2_1_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_1_2(1,1)(PERCISION) & MULTS_2_1_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(1,1)<=signed(MULTS_2_2_1(1,1)(PERCISION) & MULTS_2_2_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_2_2(1,1)(PERCISION) & MULTS_2_2_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(1,1)<=signed(MULTS_2_3_1(1,1)(PERCISION) & MULTS_2_3_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_3_2(1,1)(PERCISION) & MULTS_2_3_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(1,1)<=signed(MULTS_2_4_1(1,1)(PERCISION) & MULTS_2_4_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_4_2(1,1)(PERCISION) & MULTS_2_4_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(1,1)<=signed(MULTS_2_5_1(1,1)(PERCISION) & MULTS_2_5_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_5_2(1,1)(PERCISION) & MULTS_2_5_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(1,1)<=signed(MULTS_2_6_1(1,1)(PERCISION) & MULTS_2_6_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_6_2(1,1)(PERCISION) & MULTS_2_6_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(1,1)<=signed(MULTS_2_7_1(1,1)(PERCISION) & MULTS_2_7_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_7_2(1,1)(PERCISION) & MULTS_2_7_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(1,1)<=signed(MULTS_2_8_1(1,1)(PERCISION) & MULTS_2_8_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_8_2(1,1)(PERCISION) & MULTS_2_8_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(1,1)<=signed(MULTS_2_9_1(1,1)(PERCISION) & MULTS_2_9_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_9_2(1,1)(PERCISION) & MULTS_2_9_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(1,1)<=signed(MULTS_2_10_1(1,1)(PERCISION) & MULTS_2_10_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_10_2(1,1)(PERCISION) & MULTS_2_10_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(1,1)<=signed(MULTS_2_11_1(1,1)(PERCISION) & MULTS_2_11_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_11_2(1,1)(PERCISION) & MULTS_2_11_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(1,1)<=signed(MULTS_2_12_1(1,1)(PERCISION) & MULTS_2_12_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_12_2(1,1)(PERCISION) & MULTS_2_12_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(1,1)<=signed(MULTS_2_13_1(1,1)(PERCISION) & MULTS_2_13_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_13_2(1,1)(PERCISION) & MULTS_2_13_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(1,1)<=signed(MULTS_2_14_1(1,1)(PERCISION) & MULTS_2_14_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_14_2(1,1)(PERCISION) & MULTS_2_14_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(1,1)<=signed(MULTS_2_15_1(1,1)(PERCISION) & MULTS_2_15_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_15_2(1,1)(PERCISION) & MULTS_2_15_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(1,1)<=signed(MULTS_2_16_1(1,1)(PERCISION) & MULTS_2_16_1(1,1)(PERCISION downto 1)) + signed(MULTS_2_16_2(1,1)(PERCISION) & MULTS_2_16_2(1,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(1,1) ------------------

			MULTS_3_1_1(1,2)<=signed(MULTS_2_1_1(1,2)(PERCISION) & MULTS_2_1_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_1_2(1,2)(PERCISION) & MULTS_2_1_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(1,2)<=signed(MULTS_2_2_1(1,2)(PERCISION) & MULTS_2_2_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_2_2(1,2)(PERCISION) & MULTS_2_2_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(1,2)<=signed(MULTS_2_3_1(1,2)(PERCISION) & MULTS_2_3_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_3_2(1,2)(PERCISION) & MULTS_2_3_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(1,2)<=signed(MULTS_2_4_1(1,2)(PERCISION) & MULTS_2_4_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_4_2(1,2)(PERCISION) & MULTS_2_4_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(1,2)<=signed(MULTS_2_5_1(1,2)(PERCISION) & MULTS_2_5_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_5_2(1,2)(PERCISION) & MULTS_2_5_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(1,2)<=signed(MULTS_2_6_1(1,2)(PERCISION) & MULTS_2_6_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_6_2(1,2)(PERCISION) & MULTS_2_6_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(1,2)<=signed(MULTS_2_7_1(1,2)(PERCISION) & MULTS_2_7_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_7_2(1,2)(PERCISION) & MULTS_2_7_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(1,2)<=signed(MULTS_2_8_1(1,2)(PERCISION) & MULTS_2_8_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_8_2(1,2)(PERCISION) & MULTS_2_8_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(1,2)<=signed(MULTS_2_9_1(1,2)(PERCISION) & MULTS_2_9_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_9_2(1,2)(PERCISION) & MULTS_2_9_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(1,2)<=signed(MULTS_2_10_1(1,2)(PERCISION) & MULTS_2_10_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_10_2(1,2)(PERCISION) & MULTS_2_10_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(1,2)<=signed(MULTS_2_11_1(1,2)(PERCISION) & MULTS_2_11_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_11_2(1,2)(PERCISION) & MULTS_2_11_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(1,2)<=signed(MULTS_2_12_1(1,2)(PERCISION) & MULTS_2_12_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_12_2(1,2)(PERCISION) & MULTS_2_12_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(1,2)<=signed(MULTS_2_13_1(1,2)(PERCISION) & MULTS_2_13_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_13_2(1,2)(PERCISION) & MULTS_2_13_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(1,2)<=signed(MULTS_2_14_1(1,2)(PERCISION) & MULTS_2_14_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_14_2(1,2)(PERCISION) & MULTS_2_14_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(1,2)<=signed(MULTS_2_15_1(1,2)(PERCISION) & MULTS_2_15_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_15_2(1,2)(PERCISION) & MULTS_2_15_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(1,2)<=signed(MULTS_2_16_1(1,2)(PERCISION) & MULTS_2_16_1(1,2)(PERCISION downto 1)) + signed(MULTS_2_16_2(1,2)(PERCISION) & MULTS_2_16_2(1,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(1,2) ------------------

			MULTS_3_1_1(1,3)<=signed(MULTS_2_1_1(1,3)(PERCISION) & MULTS_2_1_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_1_2(1,3)(PERCISION) & MULTS_2_1_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(1,3)<=signed(MULTS_2_2_1(1,3)(PERCISION) & MULTS_2_2_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_2_2(1,3)(PERCISION) & MULTS_2_2_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(1,3)<=signed(MULTS_2_3_1(1,3)(PERCISION) & MULTS_2_3_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_3_2(1,3)(PERCISION) & MULTS_2_3_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(1,3)<=signed(MULTS_2_4_1(1,3)(PERCISION) & MULTS_2_4_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_4_2(1,3)(PERCISION) & MULTS_2_4_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(1,3)<=signed(MULTS_2_5_1(1,3)(PERCISION) & MULTS_2_5_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_5_2(1,3)(PERCISION) & MULTS_2_5_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(1,3)<=signed(MULTS_2_6_1(1,3)(PERCISION) & MULTS_2_6_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_6_2(1,3)(PERCISION) & MULTS_2_6_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(1,3)<=signed(MULTS_2_7_1(1,3)(PERCISION) & MULTS_2_7_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_7_2(1,3)(PERCISION) & MULTS_2_7_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(1,3)<=signed(MULTS_2_8_1(1,3)(PERCISION) & MULTS_2_8_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_8_2(1,3)(PERCISION) & MULTS_2_8_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(1,3)<=signed(MULTS_2_9_1(1,3)(PERCISION) & MULTS_2_9_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_9_2(1,3)(PERCISION) & MULTS_2_9_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(1,3)<=signed(MULTS_2_10_1(1,3)(PERCISION) & MULTS_2_10_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_10_2(1,3)(PERCISION) & MULTS_2_10_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(1,3)<=signed(MULTS_2_11_1(1,3)(PERCISION) & MULTS_2_11_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_11_2(1,3)(PERCISION) & MULTS_2_11_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(1,3)<=signed(MULTS_2_12_1(1,3)(PERCISION) & MULTS_2_12_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_12_2(1,3)(PERCISION) & MULTS_2_12_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(1,3)<=signed(MULTS_2_13_1(1,3)(PERCISION) & MULTS_2_13_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_13_2(1,3)(PERCISION) & MULTS_2_13_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(1,3)<=signed(MULTS_2_14_1(1,3)(PERCISION) & MULTS_2_14_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_14_2(1,3)(PERCISION) & MULTS_2_14_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(1,3)<=signed(MULTS_2_15_1(1,3)(PERCISION) & MULTS_2_15_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_15_2(1,3)(PERCISION) & MULTS_2_15_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(1,3)<=signed(MULTS_2_16_1(1,3)(PERCISION) & MULTS_2_16_1(1,3)(PERCISION downto 1)) + signed(MULTS_2_16_2(1,3)(PERCISION) & MULTS_2_16_2(1,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(1,3) ------------------

			MULTS_3_1_1(1,4)<=signed(MULTS_2_1_1(1,4)(PERCISION) & MULTS_2_1_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_1_2(1,4)(PERCISION) & MULTS_2_1_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(1,4)<=signed(MULTS_2_2_1(1,4)(PERCISION) & MULTS_2_2_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_2_2(1,4)(PERCISION) & MULTS_2_2_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(1,4)<=signed(MULTS_2_3_1(1,4)(PERCISION) & MULTS_2_3_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_3_2(1,4)(PERCISION) & MULTS_2_3_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(1,4)<=signed(MULTS_2_4_1(1,4)(PERCISION) & MULTS_2_4_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_4_2(1,4)(PERCISION) & MULTS_2_4_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(1,4)<=signed(MULTS_2_5_1(1,4)(PERCISION) & MULTS_2_5_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_5_2(1,4)(PERCISION) & MULTS_2_5_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(1,4)<=signed(MULTS_2_6_1(1,4)(PERCISION) & MULTS_2_6_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_6_2(1,4)(PERCISION) & MULTS_2_6_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(1,4)<=signed(MULTS_2_7_1(1,4)(PERCISION) & MULTS_2_7_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_7_2(1,4)(PERCISION) & MULTS_2_7_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(1,4)<=signed(MULTS_2_8_1(1,4)(PERCISION) & MULTS_2_8_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_8_2(1,4)(PERCISION) & MULTS_2_8_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(1,4)<=signed(MULTS_2_9_1(1,4)(PERCISION) & MULTS_2_9_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_9_2(1,4)(PERCISION) & MULTS_2_9_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(1,4)<=signed(MULTS_2_10_1(1,4)(PERCISION) & MULTS_2_10_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_10_2(1,4)(PERCISION) & MULTS_2_10_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(1,4)<=signed(MULTS_2_11_1(1,4)(PERCISION) & MULTS_2_11_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_11_2(1,4)(PERCISION) & MULTS_2_11_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(1,4)<=signed(MULTS_2_12_1(1,4)(PERCISION) & MULTS_2_12_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_12_2(1,4)(PERCISION) & MULTS_2_12_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(1,4)<=signed(MULTS_2_13_1(1,4)(PERCISION) & MULTS_2_13_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_13_2(1,4)(PERCISION) & MULTS_2_13_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(1,4)<=signed(MULTS_2_14_1(1,4)(PERCISION) & MULTS_2_14_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_14_2(1,4)(PERCISION) & MULTS_2_14_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(1,4)<=signed(MULTS_2_15_1(1,4)(PERCISION) & MULTS_2_15_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_15_2(1,4)(PERCISION) & MULTS_2_15_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(1,4)<=signed(MULTS_2_16_1(1,4)(PERCISION) & MULTS_2_16_1(1,4)(PERCISION downto 1)) + signed(MULTS_2_16_2(1,4)(PERCISION) & MULTS_2_16_2(1,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(1,4) ------------------

			MULTS_3_1_1(2,0)<=signed(MULTS_2_1_1(2,0)(PERCISION) & MULTS_2_1_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_1_2(2,0)(PERCISION) & MULTS_2_1_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(2,0)<=signed(MULTS_2_2_1(2,0)(PERCISION) & MULTS_2_2_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_2_2(2,0)(PERCISION) & MULTS_2_2_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(2,0)<=signed(MULTS_2_3_1(2,0)(PERCISION) & MULTS_2_3_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_3_2(2,0)(PERCISION) & MULTS_2_3_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(2,0)<=signed(MULTS_2_4_1(2,0)(PERCISION) & MULTS_2_4_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_4_2(2,0)(PERCISION) & MULTS_2_4_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(2,0)<=signed(MULTS_2_5_1(2,0)(PERCISION) & MULTS_2_5_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_5_2(2,0)(PERCISION) & MULTS_2_5_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(2,0)<=signed(MULTS_2_6_1(2,0)(PERCISION) & MULTS_2_6_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_6_2(2,0)(PERCISION) & MULTS_2_6_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(2,0)<=signed(MULTS_2_7_1(2,0)(PERCISION) & MULTS_2_7_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_7_2(2,0)(PERCISION) & MULTS_2_7_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(2,0)<=signed(MULTS_2_8_1(2,0)(PERCISION) & MULTS_2_8_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_8_2(2,0)(PERCISION) & MULTS_2_8_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(2,0)<=signed(MULTS_2_9_1(2,0)(PERCISION) & MULTS_2_9_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_9_2(2,0)(PERCISION) & MULTS_2_9_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(2,0)<=signed(MULTS_2_10_1(2,0)(PERCISION) & MULTS_2_10_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_10_2(2,0)(PERCISION) & MULTS_2_10_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(2,0)<=signed(MULTS_2_11_1(2,0)(PERCISION) & MULTS_2_11_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_11_2(2,0)(PERCISION) & MULTS_2_11_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(2,0)<=signed(MULTS_2_12_1(2,0)(PERCISION) & MULTS_2_12_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_12_2(2,0)(PERCISION) & MULTS_2_12_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(2,0)<=signed(MULTS_2_13_1(2,0)(PERCISION) & MULTS_2_13_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_13_2(2,0)(PERCISION) & MULTS_2_13_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(2,0)<=signed(MULTS_2_14_1(2,0)(PERCISION) & MULTS_2_14_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_14_2(2,0)(PERCISION) & MULTS_2_14_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(2,0)<=signed(MULTS_2_15_1(2,0)(PERCISION) & MULTS_2_15_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_15_2(2,0)(PERCISION) & MULTS_2_15_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(2,0)<=signed(MULTS_2_16_1(2,0)(PERCISION) & MULTS_2_16_1(2,0)(PERCISION downto 1)) + signed(MULTS_2_16_2(2,0)(PERCISION) & MULTS_2_16_2(2,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(2,0) ------------------

			MULTS_3_1_1(2,1)<=signed(MULTS_2_1_1(2,1)(PERCISION) & MULTS_2_1_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_1_2(2,1)(PERCISION) & MULTS_2_1_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(2,1)<=signed(MULTS_2_2_1(2,1)(PERCISION) & MULTS_2_2_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_2_2(2,1)(PERCISION) & MULTS_2_2_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(2,1)<=signed(MULTS_2_3_1(2,1)(PERCISION) & MULTS_2_3_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_3_2(2,1)(PERCISION) & MULTS_2_3_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(2,1)<=signed(MULTS_2_4_1(2,1)(PERCISION) & MULTS_2_4_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_4_2(2,1)(PERCISION) & MULTS_2_4_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(2,1)<=signed(MULTS_2_5_1(2,1)(PERCISION) & MULTS_2_5_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_5_2(2,1)(PERCISION) & MULTS_2_5_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(2,1)<=signed(MULTS_2_6_1(2,1)(PERCISION) & MULTS_2_6_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_6_2(2,1)(PERCISION) & MULTS_2_6_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(2,1)<=signed(MULTS_2_7_1(2,1)(PERCISION) & MULTS_2_7_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_7_2(2,1)(PERCISION) & MULTS_2_7_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(2,1)<=signed(MULTS_2_8_1(2,1)(PERCISION) & MULTS_2_8_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_8_2(2,1)(PERCISION) & MULTS_2_8_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(2,1)<=signed(MULTS_2_9_1(2,1)(PERCISION) & MULTS_2_9_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_9_2(2,1)(PERCISION) & MULTS_2_9_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(2,1)<=signed(MULTS_2_10_1(2,1)(PERCISION) & MULTS_2_10_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_10_2(2,1)(PERCISION) & MULTS_2_10_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(2,1)<=signed(MULTS_2_11_1(2,1)(PERCISION) & MULTS_2_11_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_11_2(2,1)(PERCISION) & MULTS_2_11_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(2,1)<=signed(MULTS_2_12_1(2,1)(PERCISION) & MULTS_2_12_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_12_2(2,1)(PERCISION) & MULTS_2_12_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(2,1)<=signed(MULTS_2_13_1(2,1)(PERCISION) & MULTS_2_13_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_13_2(2,1)(PERCISION) & MULTS_2_13_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(2,1)<=signed(MULTS_2_14_1(2,1)(PERCISION) & MULTS_2_14_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_14_2(2,1)(PERCISION) & MULTS_2_14_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(2,1)<=signed(MULTS_2_15_1(2,1)(PERCISION) & MULTS_2_15_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_15_2(2,1)(PERCISION) & MULTS_2_15_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(2,1)<=signed(MULTS_2_16_1(2,1)(PERCISION) & MULTS_2_16_1(2,1)(PERCISION downto 1)) + signed(MULTS_2_16_2(2,1)(PERCISION) & MULTS_2_16_2(2,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(2,1) ------------------

			MULTS_3_1_1(2,2)<=signed(MULTS_2_1_1(2,2)(PERCISION) & MULTS_2_1_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_1_2(2,2)(PERCISION) & MULTS_2_1_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(2,2)<=signed(MULTS_2_2_1(2,2)(PERCISION) & MULTS_2_2_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_2_2(2,2)(PERCISION) & MULTS_2_2_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(2,2)<=signed(MULTS_2_3_1(2,2)(PERCISION) & MULTS_2_3_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_3_2(2,2)(PERCISION) & MULTS_2_3_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(2,2)<=signed(MULTS_2_4_1(2,2)(PERCISION) & MULTS_2_4_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_4_2(2,2)(PERCISION) & MULTS_2_4_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(2,2)<=signed(MULTS_2_5_1(2,2)(PERCISION) & MULTS_2_5_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_5_2(2,2)(PERCISION) & MULTS_2_5_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(2,2)<=signed(MULTS_2_6_1(2,2)(PERCISION) & MULTS_2_6_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_6_2(2,2)(PERCISION) & MULTS_2_6_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(2,2)<=signed(MULTS_2_7_1(2,2)(PERCISION) & MULTS_2_7_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_7_2(2,2)(PERCISION) & MULTS_2_7_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(2,2)<=signed(MULTS_2_8_1(2,2)(PERCISION) & MULTS_2_8_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_8_2(2,2)(PERCISION) & MULTS_2_8_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(2,2)<=signed(MULTS_2_9_1(2,2)(PERCISION) & MULTS_2_9_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_9_2(2,2)(PERCISION) & MULTS_2_9_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(2,2)<=signed(MULTS_2_10_1(2,2)(PERCISION) & MULTS_2_10_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_10_2(2,2)(PERCISION) & MULTS_2_10_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(2,2)<=signed(MULTS_2_11_1(2,2)(PERCISION) & MULTS_2_11_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_11_2(2,2)(PERCISION) & MULTS_2_11_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(2,2)<=signed(MULTS_2_12_1(2,2)(PERCISION) & MULTS_2_12_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_12_2(2,2)(PERCISION) & MULTS_2_12_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(2,2)<=signed(MULTS_2_13_1(2,2)(PERCISION) & MULTS_2_13_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_13_2(2,2)(PERCISION) & MULTS_2_13_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(2,2)<=signed(MULTS_2_14_1(2,2)(PERCISION) & MULTS_2_14_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_14_2(2,2)(PERCISION) & MULTS_2_14_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(2,2)<=signed(MULTS_2_15_1(2,2)(PERCISION) & MULTS_2_15_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_15_2(2,2)(PERCISION) & MULTS_2_15_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(2,2)<=signed(MULTS_2_16_1(2,2)(PERCISION) & MULTS_2_16_1(2,2)(PERCISION downto 1)) + signed(MULTS_2_16_2(2,2)(PERCISION) & MULTS_2_16_2(2,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(2,2) ------------------

			MULTS_3_1_1(2,3)<=signed(MULTS_2_1_1(2,3)(PERCISION) & MULTS_2_1_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_1_2(2,3)(PERCISION) & MULTS_2_1_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(2,3)<=signed(MULTS_2_2_1(2,3)(PERCISION) & MULTS_2_2_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_2_2(2,3)(PERCISION) & MULTS_2_2_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(2,3)<=signed(MULTS_2_3_1(2,3)(PERCISION) & MULTS_2_3_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_3_2(2,3)(PERCISION) & MULTS_2_3_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(2,3)<=signed(MULTS_2_4_1(2,3)(PERCISION) & MULTS_2_4_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_4_2(2,3)(PERCISION) & MULTS_2_4_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(2,3)<=signed(MULTS_2_5_1(2,3)(PERCISION) & MULTS_2_5_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_5_2(2,3)(PERCISION) & MULTS_2_5_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(2,3)<=signed(MULTS_2_6_1(2,3)(PERCISION) & MULTS_2_6_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_6_2(2,3)(PERCISION) & MULTS_2_6_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(2,3)<=signed(MULTS_2_7_1(2,3)(PERCISION) & MULTS_2_7_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_7_2(2,3)(PERCISION) & MULTS_2_7_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(2,3)<=signed(MULTS_2_8_1(2,3)(PERCISION) & MULTS_2_8_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_8_2(2,3)(PERCISION) & MULTS_2_8_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(2,3)<=signed(MULTS_2_9_1(2,3)(PERCISION) & MULTS_2_9_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_9_2(2,3)(PERCISION) & MULTS_2_9_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(2,3)<=signed(MULTS_2_10_1(2,3)(PERCISION) & MULTS_2_10_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_10_2(2,3)(PERCISION) & MULTS_2_10_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(2,3)<=signed(MULTS_2_11_1(2,3)(PERCISION) & MULTS_2_11_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_11_2(2,3)(PERCISION) & MULTS_2_11_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(2,3)<=signed(MULTS_2_12_1(2,3)(PERCISION) & MULTS_2_12_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_12_2(2,3)(PERCISION) & MULTS_2_12_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(2,3)<=signed(MULTS_2_13_1(2,3)(PERCISION) & MULTS_2_13_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_13_2(2,3)(PERCISION) & MULTS_2_13_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(2,3)<=signed(MULTS_2_14_1(2,3)(PERCISION) & MULTS_2_14_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_14_2(2,3)(PERCISION) & MULTS_2_14_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(2,3)<=signed(MULTS_2_15_1(2,3)(PERCISION) & MULTS_2_15_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_15_2(2,3)(PERCISION) & MULTS_2_15_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(2,3)<=signed(MULTS_2_16_1(2,3)(PERCISION) & MULTS_2_16_1(2,3)(PERCISION downto 1)) + signed(MULTS_2_16_2(2,3)(PERCISION) & MULTS_2_16_2(2,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(2,3) ------------------

			MULTS_3_1_1(2,4)<=signed(MULTS_2_1_1(2,4)(PERCISION) & MULTS_2_1_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_1_2(2,4)(PERCISION) & MULTS_2_1_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(2,4)<=signed(MULTS_2_2_1(2,4)(PERCISION) & MULTS_2_2_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_2_2(2,4)(PERCISION) & MULTS_2_2_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(2,4)<=signed(MULTS_2_3_1(2,4)(PERCISION) & MULTS_2_3_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_3_2(2,4)(PERCISION) & MULTS_2_3_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(2,4)<=signed(MULTS_2_4_1(2,4)(PERCISION) & MULTS_2_4_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_4_2(2,4)(PERCISION) & MULTS_2_4_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(2,4)<=signed(MULTS_2_5_1(2,4)(PERCISION) & MULTS_2_5_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_5_2(2,4)(PERCISION) & MULTS_2_5_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(2,4)<=signed(MULTS_2_6_1(2,4)(PERCISION) & MULTS_2_6_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_6_2(2,4)(PERCISION) & MULTS_2_6_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(2,4)<=signed(MULTS_2_7_1(2,4)(PERCISION) & MULTS_2_7_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_7_2(2,4)(PERCISION) & MULTS_2_7_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(2,4)<=signed(MULTS_2_8_1(2,4)(PERCISION) & MULTS_2_8_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_8_2(2,4)(PERCISION) & MULTS_2_8_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(2,4)<=signed(MULTS_2_9_1(2,4)(PERCISION) & MULTS_2_9_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_9_2(2,4)(PERCISION) & MULTS_2_9_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(2,4)<=signed(MULTS_2_10_1(2,4)(PERCISION) & MULTS_2_10_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_10_2(2,4)(PERCISION) & MULTS_2_10_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(2,4)<=signed(MULTS_2_11_1(2,4)(PERCISION) & MULTS_2_11_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_11_2(2,4)(PERCISION) & MULTS_2_11_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(2,4)<=signed(MULTS_2_12_1(2,4)(PERCISION) & MULTS_2_12_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_12_2(2,4)(PERCISION) & MULTS_2_12_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(2,4)<=signed(MULTS_2_13_1(2,4)(PERCISION) & MULTS_2_13_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_13_2(2,4)(PERCISION) & MULTS_2_13_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(2,4)<=signed(MULTS_2_14_1(2,4)(PERCISION) & MULTS_2_14_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_14_2(2,4)(PERCISION) & MULTS_2_14_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(2,4)<=signed(MULTS_2_15_1(2,4)(PERCISION) & MULTS_2_15_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_15_2(2,4)(PERCISION) & MULTS_2_15_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(2,4)<=signed(MULTS_2_16_1(2,4)(PERCISION) & MULTS_2_16_1(2,4)(PERCISION downto 1)) + signed(MULTS_2_16_2(2,4)(PERCISION) & MULTS_2_16_2(2,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(2,4) ------------------

			MULTS_3_1_1(3,0)<=signed(MULTS_2_1_1(3,0)(PERCISION) & MULTS_2_1_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_1_2(3,0)(PERCISION) & MULTS_2_1_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(3,0)<=signed(MULTS_2_2_1(3,0)(PERCISION) & MULTS_2_2_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_2_2(3,0)(PERCISION) & MULTS_2_2_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(3,0)<=signed(MULTS_2_3_1(3,0)(PERCISION) & MULTS_2_3_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_3_2(3,0)(PERCISION) & MULTS_2_3_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(3,0)<=signed(MULTS_2_4_1(3,0)(PERCISION) & MULTS_2_4_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_4_2(3,0)(PERCISION) & MULTS_2_4_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(3,0)<=signed(MULTS_2_5_1(3,0)(PERCISION) & MULTS_2_5_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_5_2(3,0)(PERCISION) & MULTS_2_5_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(3,0)<=signed(MULTS_2_6_1(3,0)(PERCISION) & MULTS_2_6_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_6_2(3,0)(PERCISION) & MULTS_2_6_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(3,0)<=signed(MULTS_2_7_1(3,0)(PERCISION) & MULTS_2_7_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_7_2(3,0)(PERCISION) & MULTS_2_7_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(3,0)<=signed(MULTS_2_8_1(3,0)(PERCISION) & MULTS_2_8_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_8_2(3,0)(PERCISION) & MULTS_2_8_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(3,0)<=signed(MULTS_2_9_1(3,0)(PERCISION) & MULTS_2_9_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_9_2(3,0)(PERCISION) & MULTS_2_9_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(3,0)<=signed(MULTS_2_10_1(3,0)(PERCISION) & MULTS_2_10_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_10_2(3,0)(PERCISION) & MULTS_2_10_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(3,0)<=signed(MULTS_2_11_1(3,0)(PERCISION) & MULTS_2_11_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_11_2(3,0)(PERCISION) & MULTS_2_11_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(3,0)<=signed(MULTS_2_12_1(3,0)(PERCISION) & MULTS_2_12_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_12_2(3,0)(PERCISION) & MULTS_2_12_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(3,0)<=signed(MULTS_2_13_1(3,0)(PERCISION) & MULTS_2_13_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_13_2(3,0)(PERCISION) & MULTS_2_13_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(3,0)<=signed(MULTS_2_14_1(3,0)(PERCISION) & MULTS_2_14_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_14_2(3,0)(PERCISION) & MULTS_2_14_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(3,0)<=signed(MULTS_2_15_1(3,0)(PERCISION) & MULTS_2_15_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_15_2(3,0)(PERCISION) & MULTS_2_15_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(3,0)<=signed(MULTS_2_16_1(3,0)(PERCISION) & MULTS_2_16_1(3,0)(PERCISION downto 1)) + signed(MULTS_2_16_2(3,0)(PERCISION) & MULTS_2_16_2(3,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(3,0) ------------------

			MULTS_3_1_1(3,1)<=signed(MULTS_2_1_1(3,1)(PERCISION) & MULTS_2_1_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_1_2(3,1)(PERCISION) & MULTS_2_1_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(3,1)<=signed(MULTS_2_2_1(3,1)(PERCISION) & MULTS_2_2_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_2_2(3,1)(PERCISION) & MULTS_2_2_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(3,1)<=signed(MULTS_2_3_1(3,1)(PERCISION) & MULTS_2_3_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_3_2(3,1)(PERCISION) & MULTS_2_3_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(3,1)<=signed(MULTS_2_4_1(3,1)(PERCISION) & MULTS_2_4_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_4_2(3,1)(PERCISION) & MULTS_2_4_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(3,1)<=signed(MULTS_2_5_1(3,1)(PERCISION) & MULTS_2_5_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_5_2(3,1)(PERCISION) & MULTS_2_5_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(3,1)<=signed(MULTS_2_6_1(3,1)(PERCISION) & MULTS_2_6_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_6_2(3,1)(PERCISION) & MULTS_2_6_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(3,1)<=signed(MULTS_2_7_1(3,1)(PERCISION) & MULTS_2_7_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_7_2(3,1)(PERCISION) & MULTS_2_7_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(3,1)<=signed(MULTS_2_8_1(3,1)(PERCISION) & MULTS_2_8_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_8_2(3,1)(PERCISION) & MULTS_2_8_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(3,1)<=signed(MULTS_2_9_1(3,1)(PERCISION) & MULTS_2_9_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_9_2(3,1)(PERCISION) & MULTS_2_9_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(3,1)<=signed(MULTS_2_10_1(3,1)(PERCISION) & MULTS_2_10_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_10_2(3,1)(PERCISION) & MULTS_2_10_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(3,1)<=signed(MULTS_2_11_1(3,1)(PERCISION) & MULTS_2_11_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_11_2(3,1)(PERCISION) & MULTS_2_11_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(3,1)<=signed(MULTS_2_12_1(3,1)(PERCISION) & MULTS_2_12_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_12_2(3,1)(PERCISION) & MULTS_2_12_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(3,1)<=signed(MULTS_2_13_1(3,1)(PERCISION) & MULTS_2_13_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_13_2(3,1)(PERCISION) & MULTS_2_13_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(3,1)<=signed(MULTS_2_14_1(3,1)(PERCISION) & MULTS_2_14_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_14_2(3,1)(PERCISION) & MULTS_2_14_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(3,1)<=signed(MULTS_2_15_1(3,1)(PERCISION) & MULTS_2_15_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_15_2(3,1)(PERCISION) & MULTS_2_15_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(3,1)<=signed(MULTS_2_16_1(3,1)(PERCISION) & MULTS_2_16_1(3,1)(PERCISION downto 1)) + signed(MULTS_2_16_2(3,1)(PERCISION) & MULTS_2_16_2(3,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(3,1) ------------------

			MULTS_3_1_1(3,2)<=signed(MULTS_2_1_1(3,2)(PERCISION) & MULTS_2_1_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_1_2(3,2)(PERCISION) & MULTS_2_1_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(3,2)<=signed(MULTS_2_2_1(3,2)(PERCISION) & MULTS_2_2_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_2_2(3,2)(PERCISION) & MULTS_2_2_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(3,2)<=signed(MULTS_2_3_1(3,2)(PERCISION) & MULTS_2_3_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_3_2(3,2)(PERCISION) & MULTS_2_3_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(3,2)<=signed(MULTS_2_4_1(3,2)(PERCISION) & MULTS_2_4_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_4_2(3,2)(PERCISION) & MULTS_2_4_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(3,2)<=signed(MULTS_2_5_1(3,2)(PERCISION) & MULTS_2_5_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_5_2(3,2)(PERCISION) & MULTS_2_5_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(3,2)<=signed(MULTS_2_6_1(3,2)(PERCISION) & MULTS_2_6_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_6_2(3,2)(PERCISION) & MULTS_2_6_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(3,2)<=signed(MULTS_2_7_1(3,2)(PERCISION) & MULTS_2_7_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_7_2(3,2)(PERCISION) & MULTS_2_7_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(3,2)<=signed(MULTS_2_8_1(3,2)(PERCISION) & MULTS_2_8_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_8_2(3,2)(PERCISION) & MULTS_2_8_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(3,2)<=signed(MULTS_2_9_1(3,2)(PERCISION) & MULTS_2_9_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_9_2(3,2)(PERCISION) & MULTS_2_9_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(3,2)<=signed(MULTS_2_10_1(3,2)(PERCISION) & MULTS_2_10_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_10_2(3,2)(PERCISION) & MULTS_2_10_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(3,2)<=signed(MULTS_2_11_1(3,2)(PERCISION) & MULTS_2_11_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_11_2(3,2)(PERCISION) & MULTS_2_11_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(3,2)<=signed(MULTS_2_12_1(3,2)(PERCISION) & MULTS_2_12_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_12_2(3,2)(PERCISION) & MULTS_2_12_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(3,2)<=signed(MULTS_2_13_1(3,2)(PERCISION) & MULTS_2_13_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_13_2(3,2)(PERCISION) & MULTS_2_13_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(3,2)<=signed(MULTS_2_14_1(3,2)(PERCISION) & MULTS_2_14_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_14_2(3,2)(PERCISION) & MULTS_2_14_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(3,2)<=signed(MULTS_2_15_1(3,2)(PERCISION) & MULTS_2_15_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_15_2(3,2)(PERCISION) & MULTS_2_15_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(3,2)<=signed(MULTS_2_16_1(3,2)(PERCISION) & MULTS_2_16_1(3,2)(PERCISION downto 1)) + signed(MULTS_2_16_2(3,2)(PERCISION) & MULTS_2_16_2(3,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(3,2) ------------------

			MULTS_3_1_1(3,3)<=signed(MULTS_2_1_1(3,3)(PERCISION) & MULTS_2_1_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_1_2(3,3)(PERCISION) & MULTS_2_1_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(3,3)<=signed(MULTS_2_2_1(3,3)(PERCISION) & MULTS_2_2_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_2_2(3,3)(PERCISION) & MULTS_2_2_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(3,3)<=signed(MULTS_2_3_1(3,3)(PERCISION) & MULTS_2_3_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_3_2(3,3)(PERCISION) & MULTS_2_3_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(3,3)<=signed(MULTS_2_4_1(3,3)(PERCISION) & MULTS_2_4_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_4_2(3,3)(PERCISION) & MULTS_2_4_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(3,3)<=signed(MULTS_2_5_1(3,3)(PERCISION) & MULTS_2_5_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_5_2(3,3)(PERCISION) & MULTS_2_5_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(3,3)<=signed(MULTS_2_6_1(3,3)(PERCISION) & MULTS_2_6_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_6_2(3,3)(PERCISION) & MULTS_2_6_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(3,3)<=signed(MULTS_2_7_1(3,3)(PERCISION) & MULTS_2_7_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_7_2(3,3)(PERCISION) & MULTS_2_7_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(3,3)<=signed(MULTS_2_8_1(3,3)(PERCISION) & MULTS_2_8_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_8_2(3,3)(PERCISION) & MULTS_2_8_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(3,3)<=signed(MULTS_2_9_1(3,3)(PERCISION) & MULTS_2_9_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_9_2(3,3)(PERCISION) & MULTS_2_9_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(3,3)<=signed(MULTS_2_10_1(3,3)(PERCISION) & MULTS_2_10_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_10_2(3,3)(PERCISION) & MULTS_2_10_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(3,3)<=signed(MULTS_2_11_1(3,3)(PERCISION) & MULTS_2_11_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_11_2(3,3)(PERCISION) & MULTS_2_11_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(3,3)<=signed(MULTS_2_12_1(3,3)(PERCISION) & MULTS_2_12_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_12_2(3,3)(PERCISION) & MULTS_2_12_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(3,3)<=signed(MULTS_2_13_1(3,3)(PERCISION) & MULTS_2_13_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_13_2(3,3)(PERCISION) & MULTS_2_13_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(3,3)<=signed(MULTS_2_14_1(3,3)(PERCISION) & MULTS_2_14_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_14_2(3,3)(PERCISION) & MULTS_2_14_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(3,3)<=signed(MULTS_2_15_1(3,3)(PERCISION) & MULTS_2_15_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_15_2(3,3)(PERCISION) & MULTS_2_15_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(3,3)<=signed(MULTS_2_16_1(3,3)(PERCISION) & MULTS_2_16_1(3,3)(PERCISION downto 1)) + signed(MULTS_2_16_2(3,3)(PERCISION) & MULTS_2_16_2(3,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(3,3) ------------------

			MULTS_3_1_1(3,4)<=signed(MULTS_2_1_1(3,4)(PERCISION) & MULTS_2_1_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_1_2(3,4)(PERCISION) & MULTS_2_1_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(3,4)<=signed(MULTS_2_2_1(3,4)(PERCISION) & MULTS_2_2_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_2_2(3,4)(PERCISION) & MULTS_2_2_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(3,4)<=signed(MULTS_2_3_1(3,4)(PERCISION) & MULTS_2_3_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_3_2(3,4)(PERCISION) & MULTS_2_3_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(3,4)<=signed(MULTS_2_4_1(3,4)(PERCISION) & MULTS_2_4_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_4_2(3,4)(PERCISION) & MULTS_2_4_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(3,4)<=signed(MULTS_2_5_1(3,4)(PERCISION) & MULTS_2_5_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_5_2(3,4)(PERCISION) & MULTS_2_5_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(3,4)<=signed(MULTS_2_6_1(3,4)(PERCISION) & MULTS_2_6_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_6_2(3,4)(PERCISION) & MULTS_2_6_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(3,4)<=signed(MULTS_2_7_1(3,4)(PERCISION) & MULTS_2_7_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_7_2(3,4)(PERCISION) & MULTS_2_7_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(3,4)<=signed(MULTS_2_8_1(3,4)(PERCISION) & MULTS_2_8_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_8_2(3,4)(PERCISION) & MULTS_2_8_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(3,4)<=signed(MULTS_2_9_1(3,4)(PERCISION) & MULTS_2_9_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_9_2(3,4)(PERCISION) & MULTS_2_9_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(3,4)<=signed(MULTS_2_10_1(3,4)(PERCISION) & MULTS_2_10_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_10_2(3,4)(PERCISION) & MULTS_2_10_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(3,4)<=signed(MULTS_2_11_1(3,4)(PERCISION) & MULTS_2_11_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_11_2(3,4)(PERCISION) & MULTS_2_11_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(3,4)<=signed(MULTS_2_12_1(3,4)(PERCISION) & MULTS_2_12_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_12_2(3,4)(PERCISION) & MULTS_2_12_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(3,4)<=signed(MULTS_2_13_1(3,4)(PERCISION) & MULTS_2_13_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_13_2(3,4)(PERCISION) & MULTS_2_13_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(3,4)<=signed(MULTS_2_14_1(3,4)(PERCISION) & MULTS_2_14_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_14_2(3,4)(PERCISION) & MULTS_2_14_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(3,4)<=signed(MULTS_2_15_1(3,4)(PERCISION) & MULTS_2_15_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_15_2(3,4)(PERCISION) & MULTS_2_15_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(3,4)<=signed(MULTS_2_16_1(3,4)(PERCISION) & MULTS_2_16_1(3,4)(PERCISION downto 1)) + signed(MULTS_2_16_2(3,4)(PERCISION) & MULTS_2_16_2(3,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(3,4) ------------------

			MULTS_3_1_1(4,0)<=signed(MULTS_2_1_1(4,0)(PERCISION) & MULTS_2_1_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_1_2(4,0)(PERCISION) & MULTS_2_1_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(4,0)<=signed(MULTS_2_2_1(4,0)(PERCISION) & MULTS_2_2_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_2_2(4,0)(PERCISION) & MULTS_2_2_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(4,0)<=signed(MULTS_2_3_1(4,0)(PERCISION) & MULTS_2_3_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_3_2(4,0)(PERCISION) & MULTS_2_3_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(4,0)<=signed(MULTS_2_4_1(4,0)(PERCISION) & MULTS_2_4_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_4_2(4,0)(PERCISION) & MULTS_2_4_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(4,0)<=signed(MULTS_2_5_1(4,0)(PERCISION) & MULTS_2_5_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_5_2(4,0)(PERCISION) & MULTS_2_5_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(4,0)<=signed(MULTS_2_6_1(4,0)(PERCISION) & MULTS_2_6_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_6_2(4,0)(PERCISION) & MULTS_2_6_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(4,0)<=signed(MULTS_2_7_1(4,0)(PERCISION) & MULTS_2_7_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_7_2(4,0)(PERCISION) & MULTS_2_7_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(4,0)<=signed(MULTS_2_8_1(4,0)(PERCISION) & MULTS_2_8_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_8_2(4,0)(PERCISION) & MULTS_2_8_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(4,0)<=signed(MULTS_2_9_1(4,0)(PERCISION) & MULTS_2_9_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_9_2(4,0)(PERCISION) & MULTS_2_9_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(4,0)<=signed(MULTS_2_10_1(4,0)(PERCISION) & MULTS_2_10_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_10_2(4,0)(PERCISION) & MULTS_2_10_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(4,0)<=signed(MULTS_2_11_1(4,0)(PERCISION) & MULTS_2_11_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_11_2(4,0)(PERCISION) & MULTS_2_11_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(4,0)<=signed(MULTS_2_12_1(4,0)(PERCISION) & MULTS_2_12_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_12_2(4,0)(PERCISION) & MULTS_2_12_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(4,0)<=signed(MULTS_2_13_1(4,0)(PERCISION) & MULTS_2_13_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_13_2(4,0)(PERCISION) & MULTS_2_13_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(4,0)<=signed(MULTS_2_14_1(4,0)(PERCISION) & MULTS_2_14_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_14_2(4,0)(PERCISION) & MULTS_2_14_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(4,0)<=signed(MULTS_2_15_1(4,0)(PERCISION) & MULTS_2_15_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_15_2(4,0)(PERCISION) & MULTS_2_15_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(4,0)<=signed(MULTS_2_16_1(4,0)(PERCISION) & MULTS_2_16_1(4,0)(PERCISION downto 1)) + signed(MULTS_2_16_2(4,0)(PERCISION) & MULTS_2_16_2(4,0)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(4,0) ------------------

			MULTS_3_1_1(4,1)<=signed(MULTS_2_1_1(4,1)(PERCISION) & MULTS_2_1_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_1_2(4,1)(PERCISION) & MULTS_2_1_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(4,1)<=signed(MULTS_2_2_1(4,1)(PERCISION) & MULTS_2_2_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_2_2(4,1)(PERCISION) & MULTS_2_2_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(4,1)<=signed(MULTS_2_3_1(4,1)(PERCISION) & MULTS_2_3_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_3_2(4,1)(PERCISION) & MULTS_2_3_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(4,1)<=signed(MULTS_2_4_1(4,1)(PERCISION) & MULTS_2_4_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_4_2(4,1)(PERCISION) & MULTS_2_4_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(4,1)<=signed(MULTS_2_5_1(4,1)(PERCISION) & MULTS_2_5_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_5_2(4,1)(PERCISION) & MULTS_2_5_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(4,1)<=signed(MULTS_2_6_1(4,1)(PERCISION) & MULTS_2_6_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_6_2(4,1)(PERCISION) & MULTS_2_6_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(4,1)<=signed(MULTS_2_7_1(4,1)(PERCISION) & MULTS_2_7_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_7_2(4,1)(PERCISION) & MULTS_2_7_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(4,1)<=signed(MULTS_2_8_1(4,1)(PERCISION) & MULTS_2_8_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_8_2(4,1)(PERCISION) & MULTS_2_8_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(4,1)<=signed(MULTS_2_9_1(4,1)(PERCISION) & MULTS_2_9_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_9_2(4,1)(PERCISION) & MULTS_2_9_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(4,1)<=signed(MULTS_2_10_1(4,1)(PERCISION) & MULTS_2_10_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_10_2(4,1)(PERCISION) & MULTS_2_10_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(4,1)<=signed(MULTS_2_11_1(4,1)(PERCISION) & MULTS_2_11_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_11_2(4,1)(PERCISION) & MULTS_2_11_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(4,1)<=signed(MULTS_2_12_1(4,1)(PERCISION) & MULTS_2_12_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_12_2(4,1)(PERCISION) & MULTS_2_12_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(4,1)<=signed(MULTS_2_13_1(4,1)(PERCISION) & MULTS_2_13_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_13_2(4,1)(PERCISION) & MULTS_2_13_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(4,1)<=signed(MULTS_2_14_1(4,1)(PERCISION) & MULTS_2_14_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_14_2(4,1)(PERCISION) & MULTS_2_14_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(4,1)<=signed(MULTS_2_15_1(4,1)(PERCISION) & MULTS_2_15_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_15_2(4,1)(PERCISION) & MULTS_2_15_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(4,1)<=signed(MULTS_2_16_1(4,1)(PERCISION) & MULTS_2_16_1(4,1)(PERCISION downto 1)) + signed(MULTS_2_16_2(4,1)(PERCISION) & MULTS_2_16_2(4,1)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(4,1) ------------------

			MULTS_3_1_1(4,2)<=signed(MULTS_2_1_1(4,2)(PERCISION) & MULTS_2_1_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_1_2(4,2)(PERCISION) & MULTS_2_1_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(4,2)<=signed(MULTS_2_2_1(4,2)(PERCISION) & MULTS_2_2_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_2_2(4,2)(PERCISION) & MULTS_2_2_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(4,2)<=signed(MULTS_2_3_1(4,2)(PERCISION) & MULTS_2_3_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_3_2(4,2)(PERCISION) & MULTS_2_3_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(4,2)<=signed(MULTS_2_4_1(4,2)(PERCISION) & MULTS_2_4_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_4_2(4,2)(PERCISION) & MULTS_2_4_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(4,2)<=signed(MULTS_2_5_1(4,2)(PERCISION) & MULTS_2_5_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_5_2(4,2)(PERCISION) & MULTS_2_5_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(4,2)<=signed(MULTS_2_6_1(4,2)(PERCISION) & MULTS_2_6_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_6_2(4,2)(PERCISION) & MULTS_2_6_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(4,2)<=signed(MULTS_2_7_1(4,2)(PERCISION) & MULTS_2_7_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_7_2(4,2)(PERCISION) & MULTS_2_7_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(4,2)<=signed(MULTS_2_8_1(4,2)(PERCISION) & MULTS_2_8_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_8_2(4,2)(PERCISION) & MULTS_2_8_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(4,2)<=signed(MULTS_2_9_1(4,2)(PERCISION) & MULTS_2_9_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_9_2(4,2)(PERCISION) & MULTS_2_9_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(4,2)<=signed(MULTS_2_10_1(4,2)(PERCISION) & MULTS_2_10_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_10_2(4,2)(PERCISION) & MULTS_2_10_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(4,2)<=signed(MULTS_2_11_1(4,2)(PERCISION) & MULTS_2_11_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_11_2(4,2)(PERCISION) & MULTS_2_11_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(4,2)<=signed(MULTS_2_12_1(4,2)(PERCISION) & MULTS_2_12_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_12_2(4,2)(PERCISION) & MULTS_2_12_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(4,2)<=signed(MULTS_2_13_1(4,2)(PERCISION) & MULTS_2_13_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_13_2(4,2)(PERCISION) & MULTS_2_13_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(4,2)<=signed(MULTS_2_14_1(4,2)(PERCISION) & MULTS_2_14_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_14_2(4,2)(PERCISION) & MULTS_2_14_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(4,2)<=signed(MULTS_2_15_1(4,2)(PERCISION) & MULTS_2_15_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_15_2(4,2)(PERCISION) & MULTS_2_15_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(4,2)<=signed(MULTS_2_16_1(4,2)(PERCISION) & MULTS_2_16_1(4,2)(PERCISION downto 1)) + signed(MULTS_2_16_2(4,2)(PERCISION) & MULTS_2_16_2(4,2)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(4,2) ------------------

			MULTS_3_1_1(4,3)<=signed(MULTS_2_1_1(4,3)(PERCISION) & MULTS_2_1_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_1_2(4,3)(PERCISION) & MULTS_2_1_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(4,3)<=signed(MULTS_2_2_1(4,3)(PERCISION) & MULTS_2_2_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_2_2(4,3)(PERCISION) & MULTS_2_2_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(4,3)<=signed(MULTS_2_3_1(4,3)(PERCISION) & MULTS_2_3_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_3_2(4,3)(PERCISION) & MULTS_2_3_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(4,3)<=signed(MULTS_2_4_1(4,3)(PERCISION) & MULTS_2_4_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_4_2(4,3)(PERCISION) & MULTS_2_4_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(4,3)<=signed(MULTS_2_5_1(4,3)(PERCISION) & MULTS_2_5_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_5_2(4,3)(PERCISION) & MULTS_2_5_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(4,3)<=signed(MULTS_2_6_1(4,3)(PERCISION) & MULTS_2_6_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_6_2(4,3)(PERCISION) & MULTS_2_6_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(4,3)<=signed(MULTS_2_7_1(4,3)(PERCISION) & MULTS_2_7_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_7_2(4,3)(PERCISION) & MULTS_2_7_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(4,3)<=signed(MULTS_2_8_1(4,3)(PERCISION) & MULTS_2_8_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_8_2(4,3)(PERCISION) & MULTS_2_8_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(4,3)<=signed(MULTS_2_9_1(4,3)(PERCISION) & MULTS_2_9_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_9_2(4,3)(PERCISION) & MULTS_2_9_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(4,3)<=signed(MULTS_2_10_1(4,3)(PERCISION) & MULTS_2_10_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_10_2(4,3)(PERCISION) & MULTS_2_10_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(4,3)<=signed(MULTS_2_11_1(4,3)(PERCISION) & MULTS_2_11_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_11_2(4,3)(PERCISION) & MULTS_2_11_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(4,3)<=signed(MULTS_2_12_1(4,3)(PERCISION) & MULTS_2_12_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_12_2(4,3)(PERCISION) & MULTS_2_12_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(4,3)<=signed(MULTS_2_13_1(4,3)(PERCISION) & MULTS_2_13_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_13_2(4,3)(PERCISION) & MULTS_2_13_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(4,3)<=signed(MULTS_2_14_1(4,3)(PERCISION) & MULTS_2_14_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_14_2(4,3)(PERCISION) & MULTS_2_14_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(4,3)<=signed(MULTS_2_15_1(4,3)(PERCISION) & MULTS_2_15_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_15_2(4,3)(PERCISION) & MULTS_2_15_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(4,3)<=signed(MULTS_2_16_1(4,3)(PERCISION) & MULTS_2_16_1(4,3)(PERCISION downto 1)) + signed(MULTS_2_16_2(4,3)(PERCISION) & MULTS_2_16_2(4,3)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(4,3) ------------------

			MULTS_3_1_1(4,4)<=signed(MULTS_2_1_1(4,4)(PERCISION) & MULTS_2_1_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_1_2(4,4)(PERCISION) & MULTS_2_1_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(1) -----------------------

			MULTS_3_2_1(4,4)<=signed(MULTS_2_2_1(4,4)(PERCISION) & MULTS_2_2_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_2_2(4,4)(PERCISION) & MULTS_2_2_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(2) -----------------------

			MULTS_3_3_1(4,4)<=signed(MULTS_2_3_1(4,4)(PERCISION) & MULTS_2_3_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_3_2(4,4)(PERCISION) & MULTS_2_3_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(3) -----------------------

			MULTS_3_4_1(4,4)<=signed(MULTS_2_4_1(4,4)(PERCISION) & MULTS_2_4_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_4_2(4,4)(PERCISION) & MULTS_2_4_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(4) -----------------------

			MULTS_3_5_1(4,4)<=signed(MULTS_2_5_1(4,4)(PERCISION) & MULTS_2_5_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_5_2(4,4)(PERCISION) & MULTS_2_5_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(5) -----------------------

			MULTS_3_6_1(4,4)<=signed(MULTS_2_6_1(4,4)(PERCISION) & MULTS_2_6_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_6_2(4,4)(PERCISION) & MULTS_2_6_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(6) -----------------------

			MULTS_3_7_1(4,4)<=signed(MULTS_2_7_1(4,4)(PERCISION) & MULTS_2_7_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_7_2(4,4)(PERCISION) & MULTS_2_7_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(7) -----------------------

			MULTS_3_8_1(4,4)<=signed(MULTS_2_8_1(4,4)(PERCISION) & MULTS_2_8_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_8_2(4,4)(PERCISION) & MULTS_2_8_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(8) -----------------------

			MULTS_3_9_1(4,4)<=signed(MULTS_2_9_1(4,4)(PERCISION) & MULTS_2_9_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_9_2(4,4)(PERCISION) & MULTS_2_9_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(9) -----------------------

			MULTS_3_10_1(4,4)<=signed(MULTS_2_10_1(4,4)(PERCISION) & MULTS_2_10_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_10_2(4,4)(PERCISION) & MULTS_2_10_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(10) -----------------------

			MULTS_3_11_1(4,4)<=signed(MULTS_2_11_1(4,4)(PERCISION) & MULTS_2_11_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_11_2(4,4)(PERCISION) & MULTS_2_11_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(11) -----------------------

			MULTS_3_12_1(4,4)<=signed(MULTS_2_12_1(4,4)(PERCISION) & MULTS_2_12_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_12_2(4,4)(PERCISION) & MULTS_2_12_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(12) -----------------------

			MULTS_3_13_1(4,4)<=signed(MULTS_2_13_1(4,4)(PERCISION) & MULTS_2_13_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_13_2(4,4)(PERCISION) & MULTS_2_13_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(13) -----------------------

			MULTS_3_14_1(4,4)<=signed(MULTS_2_14_1(4,4)(PERCISION) & MULTS_2_14_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_14_2(4,4)(PERCISION) & MULTS_2_14_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(14) -----------------------

			MULTS_3_15_1(4,4)<=signed(MULTS_2_15_1(4,4)(PERCISION) & MULTS_2_15_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_15_2(4,4)(PERCISION) & MULTS_2_15_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(15) -----------------------

			MULTS_3_16_1(4,4)<=signed(MULTS_2_16_1(4,4)(PERCISION) & MULTS_2_16_1(4,4)(PERCISION downto 1)) + signed(MULTS_2_16_2(4,4)(PERCISION) & MULTS_2_16_2(4,4)(PERCISION downto 1));
			---------------------SUM P_MAPS of FMAP(16) -----------------------

			-----------------------END OF INDEX(4,4) ------------------



		Enable_STAGE_1<='1';
		end if;


		------------------------- Enable ADDER-TREE START -----------------------

		if Enable_STAGE_1 = '1' then
			------------------------------------STAGE-1--------------------------------------

			ADD_DEPTH_1(0,0)<=signed(MULTS_3_1_1(0,0));
			ADD_DEPTH_1(0,1)<=signed(MULTS_3_2_1(0,0));
			ADD_DEPTH_1(0,2)<=signed(MULTS_3_3_1(0,0));
			ADD_DEPTH_1(0,3)<=signed(MULTS_3_4_1(0,0));
			ADD_DEPTH_1(0,4)<=signed(MULTS_3_5_1(0,0));
			ADD_DEPTH_1(0,5)<=signed(MULTS_3_6_1(0,0));
			ADD_DEPTH_1(0,6)<=signed(MULTS_3_7_1(0,0));
			ADD_DEPTH_1(0,7)<=signed(MULTS_3_8_1(0,0));
			ADD_DEPTH_1(0,8)<=signed(MULTS_3_9_1(0,0));
			ADD_DEPTH_1(0,9)<=signed(MULTS_3_10_1(0,0));
			ADD_DEPTH_1(0,10)<=signed(MULTS_3_11_1(0,0));
			ADD_DEPTH_1(0,11)<=signed(MULTS_3_12_1(0,0));
			ADD_DEPTH_1(0,12)<=signed(MULTS_3_13_1(0,0));
			ADD_DEPTH_1(0,13)<=signed(MULTS_3_14_1(0,0));
			ADD_DEPTH_1(0,14)<=signed(MULTS_3_15_1(0,0));
			ADD_DEPTH_1(0,15)<=signed(MULTS_3_16_1(0,0));

			ADD_DEPTH_1(1,0)<=signed(MULTS_3_1_1(1,1)) + signed(MULTS_3_1_1(2,2));
			ADD_DEPTH_1(1,1)<=signed(MULTS_3_2_1(1,1)) + signed(MULTS_3_2_1(2,2));
			ADD_DEPTH_1(1,2)<=signed(MULTS_3_3_1(1,1)) + signed(MULTS_3_3_1(2,2));
			ADD_DEPTH_1(1,3)<=signed(MULTS_3_4_1(1,1)) + signed(MULTS_3_4_1(2,2));
			ADD_DEPTH_1(1,4)<=signed(MULTS_3_5_1(1,1)) + signed(MULTS_3_5_1(2,2));
			ADD_DEPTH_1(1,5)<=signed(MULTS_3_6_1(1,1)) + signed(MULTS_3_6_1(2,2));
			ADD_DEPTH_1(1,6)<=signed(MULTS_3_7_1(1,1)) + signed(MULTS_3_7_1(2,2));
			ADD_DEPTH_1(1,7)<=signed(MULTS_3_8_1(1,1)) + signed(MULTS_3_8_1(2,2));
			ADD_DEPTH_1(1,8)<=signed(MULTS_3_9_1(1,1)) + signed(MULTS_3_9_1(2,2));
			ADD_DEPTH_1(1,9)<=signed(MULTS_3_10_1(1,1)) + signed(MULTS_3_10_1(2,2));
			ADD_DEPTH_1(1,10)<=signed(MULTS_3_11_1(1,1)) + signed(MULTS_3_11_1(2,2));
			ADD_DEPTH_1(1,11)<=signed(MULTS_3_12_1(1,1)) + signed(MULTS_3_12_1(2,2));
			ADD_DEPTH_1(1,12)<=signed(MULTS_3_13_1(1,1)) + signed(MULTS_3_13_1(2,2));
			ADD_DEPTH_1(1,13)<=signed(MULTS_3_14_1(1,1)) + signed(MULTS_3_14_1(2,2));
			ADD_DEPTH_1(1,14)<=signed(MULTS_3_15_1(1,1)) + signed(MULTS_3_15_1(2,2));
			ADD_DEPTH_1(1,15)<=signed(MULTS_3_16_1(1,1)) + signed(MULTS_3_16_1(2,2));

			ADD_DEPTH_1(2,0)<=signed(MULTS_3_1_1(3,3)) + signed(MULTS_3_1_1(4,4));
			ADD_DEPTH_1(2,1)<=signed(MULTS_3_2_1(3,3)) + signed(MULTS_3_2_1(4,4));
			ADD_DEPTH_1(2,2)<=signed(MULTS_3_3_1(3,3)) + signed(MULTS_3_3_1(4,4));
			ADD_DEPTH_1(2,3)<=signed(MULTS_3_4_1(3,3)) + signed(MULTS_3_4_1(4,4));
			ADD_DEPTH_1(2,4)<=signed(MULTS_3_5_1(3,3)) + signed(MULTS_3_5_1(4,4));
			ADD_DEPTH_1(2,5)<=signed(MULTS_3_6_1(3,3)) + signed(MULTS_3_6_1(4,4));
			ADD_DEPTH_1(2,6)<=signed(MULTS_3_7_1(3,3)) + signed(MULTS_3_7_1(4,4));
			ADD_DEPTH_1(2,7)<=signed(MULTS_3_8_1(3,3)) + signed(MULTS_3_8_1(4,4));
			ADD_DEPTH_1(2,8)<=signed(MULTS_3_9_1(3,3)) + signed(MULTS_3_9_1(4,4));
			ADD_DEPTH_1(2,9)<=signed(MULTS_3_10_1(3,3)) + signed(MULTS_3_10_1(4,4));
			ADD_DEPTH_1(2,10)<=signed(MULTS_3_11_1(3,3)) + signed(MULTS_3_11_1(4,4));
			ADD_DEPTH_1(2,11)<=signed(MULTS_3_12_1(3,3)) + signed(MULTS_3_12_1(4,4));
			ADD_DEPTH_1(2,12)<=signed(MULTS_3_13_1(3,3)) + signed(MULTS_3_13_1(4,4));
			ADD_DEPTH_1(2,13)<=signed(MULTS_3_14_1(3,3)) + signed(MULTS_3_14_1(4,4));
			ADD_DEPTH_1(2,14)<=signed(MULTS_3_15_1(3,3)) + signed(MULTS_3_15_1(4,4));
			ADD_DEPTH_1(2,15)<=signed(MULTS_3_16_1(3,3)) + signed(MULTS_3_16_1(4,4));


			ADD_DEPTH_1(3,0)<=signed(MULTS_3_1_1(0,1)) + signed(MULTS_3_1_1(1,0));
			ADD_DEPTH_1(3,1)<=signed(MULTS_3_2_1(0,1)) + signed(MULTS_3_2_1(1,0));
			ADD_DEPTH_1(3,2)<=signed(MULTS_3_3_1(0,1)) + signed(MULTS_3_3_1(1,0));
			ADD_DEPTH_1(3,3)<=signed(MULTS_3_4_1(0,1)) + signed(MULTS_3_4_1(1,0));
			ADD_DEPTH_1(3,4)<=signed(MULTS_3_5_1(0,1)) + signed(MULTS_3_5_1(1,0));
			ADD_DEPTH_1(3,5)<=signed(MULTS_3_6_1(0,1)) + signed(MULTS_3_6_1(1,0));
			ADD_DEPTH_1(3,6)<=signed(MULTS_3_7_1(0,1)) + signed(MULTS_3_7_1(1,0));
			ADD_DEPTH_1(3,7)<=signed(MULTS_3_8_1(0,1)) + signed(MULTS_3_8_1(1,0));
			ADD_DEPTH_1(3,8)<=signed(MULTS_3_9_1(0,1)) + signed(MULTS_3_9_1(1,0));
			ADD_DEPTH_1(3,9)<=signed(MULTS_3_10_1(0,1)) + signed(MULTS_3_10_1(1,0));
			ADD_DEPTH_1(3,10)<=signed(MULTS_3_11_1(0,1)) + signed(MULTS_3_11_1(1,0));
			ADD_DEPTH_1(3,11)<=signed(MULTS_3_12_1(0,1)) + signed(MULTS_3_12_1(1,0));
			ADD_DEPTH_1(3,12)<=signed(MULTS_3_13_1(0,1)) + signed(MULTS_3_13_1(1,0));
			ADD_DEPTH_1(3,13)<=signed(MULTS_3_14_1(0,1)) + signed(MULTS_3_14_1(1,0));
			ADD_DEPTH_1(3,14)<=signed(MULTS_3_15_1(0,1)) + signed(MULTS_3_15_1(1,0));
			ADD_DEPTH_1(3,15)<=signed(MULTS_3_16_1(0,1)) + signed(MULTS_3_16_1(1,0));

			ADD_DEPTH_1(4,0)<=signed(MULTS_3_1_1(0,2)) + signed(MULTS_3_1_1(2,0));
			ADD_DEPTH_1(4,1)<=signed(MULTS_3_2_1(0,2)) + signed(MULTS_3_2_1(2,0));
			ADD_DEPTH_1(4,2)<=signed(MULTS_3_3_1(0,2)) + signed(MULTS_3_3_1(2,0));
			ADD_DEPTH_1(4,3)<=signed(MULTS_3_4_1(0,2)) + signed(MULTS_3_4_1(2,0));
			ADD_DEPTH_1(4,4)<=signed(MULTS_3_5_1(0,2)) + signed(MULTS_3_5_1(2,0));
			ADD_DEPTH_1(4,5)<=signed(MULTS_3_6_1(0,2)) + signed(MULTS_3_6_1(2,0));
			ADD_DEPTH_1(4,6)<=signed(MULTS_3_7_1(0,2)) + signed(MULTS_3_7_1(2,0));
			ADD_DEPTH_1(4,7)<=signed(MULTS_3_8_1(0,2)) + signed(MULTS_3_8_1(2,0));
			ADD_DEPTH_1(4,8)<=signed(MULTS_3_9_1(0,2)) + signed(MULTS_3_9_1(2,0));
			ADD_DEPTH_1(4,9)<=signed(MULTS_3_10_1(0,2)) + signed(MULTS_3_10_1(2,0));
			ADD_DEPTH_1(4,10)<=signed(MULTS_3_11_1(0,2)) + signed(MULTS_3_11_1(2,0));
			ADD_DEPTH_1(4,11)<=signed(MULTS_3_12_1(0,2)) + signed(MULTS_3_12_1(2,0));
			ADD_DEPTH_1(4,12)<=signed(MULTS_3_13_1(0,2)) + signed(MULTS_3_13_1(2,0));
			ADD_DEPTH_1(4,13)<=signed(MULTS_3_14_1(0,2)) + signed(MULTS_3_14_1(2,0));
			ADD_DEPTH_1(4,14)<=signed(MULTS_3_15_1(0,2)) + signed(MULTS_3_15_1(2,0));
			ADD_DEPTH_1(4,15)<=signed(MULTS_3_16_1(0,2)) + signed(MULTS_3_16_1(2,0));

			ADD_DEPTH_1(5,0)<=signed(MULTS_3_1_1(0,3)) + signed(MULTS_3_1_1(3,0));
			ADD_DEPTH_1(5,1)<=signed(MULTS_3_2_1(0,3)) + signed(MULTS_3_2_1(3,0));
			ADD_DEPTH_1(5,2)<=signed(MULTS_3_3_1(0,3)) + signed(MULTS_3_3_1(3,0));
			ADD_DEPTH_1(5,3)<=signed(MULTS_3_4_1(0,3)) + signed(MULTS_3_4_1(3,0));
			ADD_DEPTH_1(5,4)<=signed(MULTS_3_5_1(0,3)) + signed(MULTS_3_5_1(3,0));
			ADD_DEPTH_1(5,5)<=signed(MULTS_3_6_1(0,3)) + signed(MULTS_3_6_1(3,0));
			ADD_DEPTH_1(5,6)<=signed(MULTS_3_7_1(0,3)) + signed(MULTS_3_7_1(3,0));
			ADD_DEPTH_1(5,7)<=signed(MULTS_3_8_1(0,3)) + signed(MULTS_3_8_1(3,0));
			ADD_DEPTH_1(5,8)<=signed(MULTS_3_9_1(0,3)) + signed(MULTS_3_9_1(3,0));
			ADD_DEPTH_1(5,9)<=signed(MULTS_3_10_1(0,3)) + signed(MULTS_3_10_1(3,0));
			ADD_DEPTH_1(5,10)<=signed(MULTS_3_11_1(0,3)) + signed(MULTS_3_11_1(3,0));
			ADD_DEPTH_1(5,11)<=signed(MULTS_3_12_1(0,3)) + signed(MULTS_3_12_1(3,0));
			ADD_DEPTH_1(5,12)<=signed(MULTS_3_13_1(0,3)) + signed(MULTS_3_13_1(3,0));
			ADD_DEPTH_1(5,13)<=signed(MULTS_3_14_1(0,3)) + signed(MULTS_3_14_1(3,0));
			ADD_DEPTH_1(5,14)<=signed(MULTS_3_15_1(0,3)) + signed(MULTS_3_15_1(3,0));
			ADD_DEPTH_1(5,15)<=signed(MULTS_3_16_1(0,3)) + signed(MULTS_3_16_1(3,0));

			ADD_DEPTH_1(6,0)<=signed(MULTS_3_1_1(0,4)) + signed(MULTS_3_1_1(4,0));
			ADD_DEPTH_1(6,1)<=signed(MULTS_3_2_1(0,4)) + signed(MULTS_3_2_1(4,0));
			ADD_DEPTH_1(6,2)<=signed(MULTS_3_3_1(0,4)) + signed(MULTS_3_3_1(4,0));
			ADD_DEPTH_1(6,3)<=signed(MULTS_3_4_1(0,4)) + signed(MULTS_3_4_1(4,0));
			ADD_DEPTH_1(6,4)<=signed(MULTS_3_5_1(0,4)) + signed(MULTS_3_5_1(4,0));
			ADD_DEPTH_1(6,5)<=signed(MULTS_3_6_1(0,4)) + signed(MULTS_3_6_1(4,0));
			ADD_DEPTH_1(6,6)<=signed(MULTS_3_7_1(0,4)) + signed(MULTS_3_7_1(4,0));
			ADD_DEPTH_1(6,7)<=signed(MULTS_3_8_1(0,4)) + signed(MULTS_3_8_1(4,0));
			ADD_DEPTH_1(6,8)<=signed(MULTS_3_9_1(0,4)) + signed(MULTS_3_9_1(4,0));
			ADD_DEPTH_1(6,9)<=signed(MULTS_3_10_1(0,4)) + signed(MULTS_3_10_1(4,0));
			ADD_DEPTH_1(6,10)<=signed(MULTS_3_11_1(0,4)) + signed(MULTS_3_11_1(4,0));
			ADD_DEPTH_1(6,11)<=signed(MULTS_3_12_1(0,4)) + signed(MULTS_3_12_1(4,0));
			ADD_DEPTH_1(6,12)<=signed(MULTS_3_13_1(0,4)) + signed(MULTS_3_13_1(4,0));
			ADD_DEPTH_1(6,13)<=signed(MULTS_3_14_1(0,4)) + signed(MULTS_3_14_1(4,0));
			ADD_DEPTH_1(6,14)<=signed(MULTS_3_15_1(0,4)) + signed(MULTS_3_15_1(4,0));
			ADD_DEPTH_1(6,15)<=signed(MULTS_3_16_1(0,4)) + signed(MULTS_3_16_1(4,0));

			ADD_DEPTH_1(7,0)<=signed(MULTS_3_1_1(1,2)) + signed(MULTS_3_1_1(2,1));
			ADD_DEPTH_1(7,1)<=signed(MULTS_3_2_1(1,2)) + signed(MULTS_3_2_1(2,1));
			ADD_DEPTH_1(7,2)<=signed(MULTS_3_3_1(1,2)) + signed(MULTS_3_3_1(2,1));
			ADD_DEPTH_1(7,3)<=signed(MULTS_3_4_1(1,2)) + signed(MULTS_3_4_1(2,1));
			ADD_DEPTH_1(7,4)<=signed(MULTS_3_5_1(1,2)) + signed(MULTS_3_5_1(2,1));
			ADD_DEPTH_1(7,5)<=signed(MULTS_3_6_1(1,2)) + signed(MULTS_3_6_1(2,1));
			ADD_DEPTH_1(7,6)<=signed(MULTS_3_7_1(1,2)) + signed(MULTS_3_7_1(2,1));
			ADD_DEPTH_1(7,7)<=signed(MULTS_3_8_1(1,2)) + signed(MULTS_3_8_1(2,1));
			ADD_DEPTH_1(7,8)<=signed(MULTS_3_9_1(1,2)) + signed(MULTS_3_9_1(2,1));
			ADD_DEPTH_1(7,9)<=signed(MULTS_3_10_1(1,2)) + signed(MULTS_3_10_1(2,1));
			ADD_DEPTH_1(7,10)<=signed(MULTS_3_11_1(1,2)) + signed(MULTS_3_11_1(2,1));
			ADD_DEPTH_1(7,11)<=signed(MULTS_3_12_1(1,2)) + signed(MULTS_3_12_1(2,1));
			ADD_DEPTH_1(7,12)<=signed(MULTS_3_13_1(1,2)) + signed(MULTS_3_13_1(2,1));
			ADD_DEPTH_1(7,13)<=signed(MULTS_3_14_1(1,2)) + signed(MULTS_3_14_1(2,1));
			ADD_DEPTH_1(7,14)<=signed(MULTS_3_15_1(1,2)) + signed(MULTS_3_15_1(2,1));
			ADD_DEPTH_1(7,15)<=signed(MULTS_3_16_1(1,2)) + signed(MULTS_3_16_1(2,1));

			ADD_DEPTH_1(8,0)<=signed(MULTS_3_1_1(1,3)) + signed(MULTS_3_1_1(3,1));
			ADD_DEPTH_1(8,1)<=signed(MULTS_3_2_1(1,3)) + signed(MULTS_3_2_1(3,1));
			ADD_DEPTH_1(8,2)<=signed(MULTS_3_3_1(1,3)) + signed(MULTS_3_3_1(3,1));
			ADD_DEPTH_1(8,3)<=signed(MULTS_3_4_1(1,3)) + signed(MULTS_3_4_1(3,1));
			ADD_DEPTH_1(8,4)<=signed(MULTS_3_5_1(1,3)) + signed(MULTS_3_5_1(3,1));
			ADD_DEPTH_1(8,5)<=signed(MULTS_3_6_1(1,3)) + signed(MULTS_3_6_1(3,1));
			ADD_DEPTH_1(8,6)<=signed(MULTS_3_7_1(1,3)) + signed(MULTS_3_7_1(3,1));
			ADD_DEPTH_1(8,7)<=signed(MULTS_3_8_1(1,3)) + signed(MULTS_3_8_1(3,1));
			ADD_DEPTH_1(8,8)<=signed(MULTS_3_9_1(1,3)) + signed(MULTS_3_9_1(3,1));
			ADD_DEPTH_1(8,9)<=signed(MULTS_3_10_1(1,3)) + signed(MULTS_3_10_1(3,1));
			ADD_DEPTH_1(8,10)<=signed(MULTS_3_11_1(1,3)) + signed(MULTS_3_11_1(3,1));
			ADD_DEPTH_1(8,11)<=signed(MULTS_3_12_1(1,3)) + signed(MULTS_3_12_1(3,1));
			ADD_DEPTH_1(8,12)<=signed(MULTS_3_13_1(1,3)) + signed(MULTS_3_13_1(3,1));
			ADD_DEPTH_1(8,13)<=signed(MULTS_3_14_1(1,3)) + signed(MULTS_3_14_1(3,1));
			ADD_DEPTH_1(8,14)<=signed(MULTS_3_15_1(1,3)) + signed(MULTS_3_15_1(3,1));
			ADD_DEPTH_1(8,15)<=signed(MULTS_3_16_1(1,3)) + signed(MULTS_3_16_1(3,1));

			ADD_DEPTH_1(9,0)<=signed(MULTS_3_1_1(1,4)) + signed(MULTS_3_1_1(4,1));
			ADD_DEPTH_1(9,1)<=signed(MULTS_3_2_1(1,4)) + signed(MULTS_3_2_1(4,1));
			ADD_DEPTH_1(9,2)<=signed(MULTS_3_3_1(1,4)) + signed(MULTS_3_3_1(4,1));
			ADD_DEPTH_1(9,3)<=signed(MULTS_3_4_1(1,4)) + signed(MULTS_3_4_1(4,1));
			ADD_DEPTH_1(9,4)<=signed(MULTS_3_5_1(1,4)) + signed(MULTS_3_5_1(4,1));
			ADD_DEPTH_1(9,5)<=signed(MULTS_3_6_1(1,4)) + signed(MULTS_3_6_1(4,1));
			ADD_DEPTH_1(9,6)<=signed(MULTS_3_7_1(1,4)) + signed(MULTS_3_7_1(4,1));
			ADD_DEPTH_1(9,7)<=signed(MULTS_3_8_1(1,4)) + signed(MULTS_3_8_1(4,1));
			ADD_DEPTH_1(9,8)<=signed(MULTS_3_9_1(1,4)) + signed(MULTS_3_9_1(4,1));
			ADD_DEPTH_1(9,9)<=signed(MULTS_3_10_1(1,4)) + signed(MULTS_3_10_1(4,1));
			ADD_DEPTH_1(9,10)<=signed(MULTS_3_11_1(1,4)) + signed(MULTS_3_11_1(4,1));
			ADD_DEPTH_1(9,11)<=signed(MULTS_3_12_1(1,4)) + signed(MULTS_3_12_1(4,1));
			ADD_DEPTH_1(9,12)<=signed(MULTS_3_13_1(1,4)) + signed(MULTS_3_13_1(4,1));
			ADD_DEPTH_1(9,13)<=signed(MULTS_3_14_1(1,4)) + signed(MULTS_3_14_1(4,1));
			ADD_DEPTH_1(9,14)<=signed(MULTS_3_15_1(1,4)) + signed(MULTS_3_15_1(4,1));
			ADD_DEPTH_1(9,15)<=signed(MULTS_3_16_1(1,4)) + signed(MULTS_3_16_1(4,1));

			ADD_DEPTH_1(10,0)<=signed(MULTS_3_1_1(2,3)) + signed(MULTS_3_1_1(3,2));
			ADD_DEPTH_1(10,1)<=signed(MULTS_3_2_1(2,3)) + signed(MULTS_3_2_1(3,2));
			ADD_DEPTH_1(10,2)<=signed(MULTS_3_3_1(2,3)) + signed(MULTS_3_3_1(3,2));
			ADD_DEPTH_1(10,3)<=signed(MULTS_3_4_1(2,3)) + signed(MULTS_3_4_1(3,2));
			ADD_DEPTH_1(10,4)<=signed(MULTS_3_5_1(2,3)) + signed(MULTS_3_5_1(3,2));
			ADD_DEPTH_1(10,5)<=signed(MULTS_3_6_1(2,3)) + signed(MULTS_3_6_1(3,2));
			ADD_DEPTH_1(10,6)<=signed(MULTS_3_7_1(2,3)) + signed(MULTS_3_7_1(3,2));
			ADD_DEPTH_1(10,7)<=signed(MULTS_3_8_1(2,3)) + signed(MULTS_3_8_1(3,2));
			ADD_DEPTH_1(10,8)<=signed(MULTS_3_9_1(2,3)) + signed(MULTS_3_9_1(3,2));
			ADD_DEPTH_1(10,9)<=signed(MULTS_3_10_1(2,3)) + signed(MULTS_3_10_1(3,2));
			ADD_DEPTH_1(10,10)<=signed(MULTS_3_11_1(2,3)) + signed(MULTS_3_11_1(3,2));
			ADD_DEPTH_1(10,11)<=signed(MULTS_3_12_1(2,3)) + signed(MULTS_3_12_1(3,2));
			ADD_DEPTH_1(10,12)<=signed(MULTS_3_13_1(2,3)) + signed(MULTS_3_13_1(3,2));
			ADD_DEPTH_1(10,13)<=signed(MULTS_3_14_1(2,3)) + signed(MULTS_3_14_1(3,2));
			ADD_DEPTH_1(10,14)<=signed(MULTS_3_15_1(2,3)) + signed(MULTS_3_15_1(3,2));
			ADD_DEPTH_1(10,15)<=signed(MULTS_3_16_1(2,3)) + signed(MULTS_3_16_1(3,2));

			ADD_DEPTH_1(11,0)<=signed(MULTS_3_1_1(2,4)) + signed(MULTS_3_1_1(4,2));
			ADD_DEPTH_1(11,1)<=signed(MULTS_3_2_1(2,4)) + signed(MULTS_3_2_1(4,2));
			ADD_DEPTH_1(11,2)<=signed(MULTS_3_3_1(2,4)) + signed(MULTS_3_3_1(4,2));
			ADD_DEPTH_1(11,3)<=signed(MULTS_3_4_1(2,4)) + signed(MULTS_3_4_1(4,2));
			ADD_DEPTH_1(11,4)<=signed(MULTS_3_5_1(2,4)) + signed(MULTS_3_5_1(4,2));
			ADD_DEPTH_1(11,5)<=signed(MULTS_3_6_1(2,4)) + signed(MULTS_3_6_1(4,2));
			ADD_DEPTH_1(11,6)<=signed(MULTS_3_7_1(2,4)) + signed(MULTS_3_7_1(4,2));
			ADD_DEPTH_1(11,7)<=signed(MULTS_3_8_1(2,4)) + signed(MULTS_3_8_1(4,2));
			ADD_DEPTH_1(11,8)<=signed(MULTS_3_9_1(2,4)) + signed(MULTS_3_9_1(4,2));
			ADD_DEPTH_1(11,9)<=signed(MULTS_3_10_1(2,4)) + signed(MULTS_3_10_1(4,2));
			ADD_DEPTH_1(11,10)<=signed(MULTS_3_11_1(2,4)) + signed(MULTS_3_11_1(4,2));
			ADD_DEPTH_1(11,11)<=signed(MULTS_3_12_1(2,4)) + signed(MULTS_3_12_1(4,2));
			ADD_DEPTH_1(11,12)<=signed(MULTS_3_13_1(2,4)) + signed(MULTS_3_13_1(4,2));
			ADD_DEPTH_1(11,13)<=signed(MULTS_3_14_1(2,4)) + signed(MULTS_3_14_1(4,2));
			ADD_DEPTH_1(11,14)<=signed(MULTS_3_15_1(2,4)) + signed(MULTS_3_15_1(4,2));
			ADD_DEPTH_1(11,15)<=signed(MULTS_3_16_1(2,4)) + signed(MULTS_3_16_1(4,2));

			ADD_DEPTH_1(12,0)<=signed(MULTS_3_1_1(3,4)) + signed(MULTS_3_1_1(4,3));
			ADD_DEPTH_1(12,1)<=signed(MULTS_3_2_1(3,4)) + signed(MULTS_3_2_1(4,3));
			ADD_DEPTH_1(12,2)<=signed(MULTS_3_3_1(3,4)) + signed(MULTS_3_3_1(4,3));
			ADD_DEPTH_1(12,3)<=signed(MULTS_3_4_1(3,4)) + signed(MULTS_3_4_1(4,3));
			ADD_DEPTH_1(12,4)<=signed(MULTS_3_5_1(3,4)) + signed(MULTS_3_5_1(4,3));
			ADD_DEPTH_1(12,5)<=signed(MULTS_3_6_1(3,4)) + signed(MULTS_3_6_1(4,3));
			ADD_DEPTH_1(12,6)<=signed(MULTS_3_7_1(3,4)) + signed(MULTS_3_7_1(4,3));
			ADD_DEPTH_1(12,7)<=signed(MULTS_3_8_1(3,4)) + signed(MULTS_3_8_1(4,3));
			ADD_DEPTH_1(12,8)<=signed(MULTS_3_9_1(3,4)) + signed(MULTS_3_9_1(4,3));
			ADD_DEPTH_1(12,9)<=signed(MULTS_3_10_1(3,4)) + signed(MULTS_3_10_1(4,3));
			ADD_DEPTH_1(12,10)<=signed(MULTS_3_11_1(3,4)) + signed(MULTS_3_11_1(4,3));
			ADD_DEPTH_1(12,11)<=signed(MULTS_3_12_1(3,4)) + signed(MULTS_3_12_1(4,3));
			ADD_DEPTH_1(12,12)<=signed(MULTS_3_13_1(3,4)) + signed(MULTS_3_13_1(4,3));
			ADD_DEPTH_1(12,13)<=signed(MULTS_3_14_1(3,4)) + signed(MULTS_3_14_1(4,3));
			ADD_DEPTH_1(12,14)<=signed(MULTS_3_15_1(3,4)) + signed(MULTS_3_15_1(4,3));
			ADD_DEPTH_1(12,15)<=signed(MULTS_3_16_1(3,4)) + signed(MULTS_3_16_1(4,3));



				Enable_STAGE_2<= '1';
			end if; 
			------------------------------------STAGE-2--------------------------------------
		if Enable_STAGE_2 = '1' then

			ADD_DEPTH_2(0,0)<=signed(ADD_DEPTH_1(0,0));
			ADD_DEPTH_2(0,1)<=signed(ADD_DEPTH_1(0,1));
			ADD_DEPTH_2(0,2)<=signed(ADD_DEPTH_1(0,2));
			ADD_DEPTH_2(0,3)<=signed(ADD_DEPTH_1(0,3));
			ADD_DEPTH_2(0,4)<=signed(ADD_DEPTH_1(0,4));
			ADD_DEPTH_2(0,5)<=signed(ADD_DEPTH_1(0,5));
			ADD_DEPTH_2(0,6)<=signed(ADD_DEPTH_1(0,6));
			ADD_DEPTH_2(0,7)<=signed(ADD_DEPTH_1(0,7));
			ADD_DEPTH_2(0,8)<=signed(ADD_DEPTH_1(0,8));
			ADD_DEPTH_2(0,9)<=signed(ADD_DEPTH_1(0,9));
			ADD_DEPTH_2(0,10)<=signed(ADD_DEPTH_1(0,10));
			ADD_DEPTH_2(0,11)<=signed(ADD_DEPTH_1(0,11));
			ADD_DEPTH_2(0,12)<=signed(ADD_DEPTH_1(0,12));
			ADD_DEPTH_2(0,13)<=signed(ADD_DEPTH_1(0,13));
			ADD_DEPTH_2(0,14)<=signed(ADD_DEPTH_1(0,14));
			ADD_DEPTH_2(0,15)<=signed(ADD_DEPTH_1(0,15));

			ADD_DEPTH_2(1,0)<=signed(ADD_DEPTH_1(1,0)) + signed(ADD_DEPTH_1(2,0));
			ADD_DEPTH_2(1,1)<=signed(ADD_DEPTH_1(1,1)) + signed(ADD_DEPTH_1(2,1));
			ADD_DEPTH_2(1,2)<=signed(ADD_DEPTH_1(1,2)) + signed(ADD_DEPTH_1(2,2));
			ADD_DEPTH_2(1,3)<=signed(ADD_DEPTH_1(1,3)) + signed(ADD_DEPTH_1(2,3));
			ADD_DEPTH_2(1,4)<=signed(ADD_DEPTH_1(1,4)) + signed(ADD_DEPTH_1(2,4));
			ADD_DEPTH_2(1,5)<=signed(ADD_DEPTH_1(1,5)) + signed(ADD_DEPTH_1(2,5));
			ADD_DEPTH_2(1,6)<=signed(ADD_DEPTH_1(1,6)) + signed(ADD_DEPTH_1(2,6));
			ADD_DEPTH_2(1,7)<=signed(ADD_DEPTH_1(1,7)) + signed(ADD_DEPTH_1(2,7));
			ADD_DEPTH_2(1,8)<=signed(ADD_DEPTH_1(1,8)) + signed(ADD_DEPTH_1(2,8));
			ADD_DEPTH_2(1,9)<=signed(ADD_DEPTH_1(1,9)) + signed(ADD_DEPTH_1(2,9));
			ADD_DEPTH_2(1,10)<=signed(ADD_DEPTH_1(1,10)) + signed(ADD_DEPTH_1(2,10));
			ADD_DEPTH_2(1,11)<=signed(ADD_DEPTH_1(1,11)) + signed(ADD_DEPTH_1(2,11));
			ADD_DEPTH_2(1,12)<=signed(ADD_DEPTH_1(1,12)) + signed(ADD_DEPTH_1(2,12));
			ADD_DEPTH_2(1,13)<=signed(ADD_DEPTH_1(1,13)) + signed(ADD_DEPTH_1(2,13));
			ADD_DEPTH_2(1,14)<=signed(ADD_DEPTH_1(1,14)) + signed(ADD_DEPTH_1(2,14));
			ADD_DEPTH_2(1,15)<=signed(ADD_DEPTH_1(1,15)) + signed(ADD_DEPTH_1(2,15));

			ADD_DEPTH_2(2,0)<=signed(ADD_DEPTH_1(3,0)) + signed(ADD_DEPTH_1(4,0));
			ADD_DEPTH_2(2,1)<=signed(ADD_DEPTH_1(3,1)) + signed(ADD_DEPTH_1(4,1));
			ADD_DEPTH_2(2,2)<=signed(ADD_DEPTH_1(3,2)) + signed(ADD_DEPTH_1(4,2));
			ADD_DEPTH_2(2,3)<=signed(ADD_DEPTH_1(3,3)) + signed(ADD_DEPTH_1(4,3));
			ADD_DEPTH_2(2,4)<=signed(ADD_DEPTH_1(3,4)) + signed(ADD_DEPTH_1(4,4));
			ADD_DEPTH_2(2,5)<=signed(ADD_DEPTH_1(3,5)) + signed(ADD_DEPTH_1(4,5));
			ADD_DEPTH_2(2,6)<=signed(ADD_DEPTH_1(3,6)) + signed(ADD_DEPTH_1(4,6));
			ADD_DEPTH_2(2,7)<=signed(ADD_DEPTH_1(3,7)) + signed(ADD_DEPTH_1(4,7));
			ADD_DEPTH_2(2,8)<=signed(ADD_DEPTH_1(3,8)) + signed(ADD_DEPTH_1(4,8));
			ADD_DEPTH_2(2,9)<=signed(ADD_DEPTH_1(3,9)) + signed(ADD_DEPTH_1(4,9));
			ADD_DEPTH_2(2,10)<=signed(ADD_DEPTH_1(3,10)) + signed(ADD_DEPTH_1(4,10));
			ADD_DEPTH_2(2,11)<=signed(ADD_DEPTH_1(3,11)) + signed(ADD_DEPTH_1(4,11));
			ADD_DEPTH_2(2,12)<=signed(ADD_DEPTH_1(3,12)) + signed(ADD_DEPTH_1(4,12));
			ADD_DEPTH_2(2,13)<=signed(ADD_DEPTH_1(3,13)) + signed(ADD_DEPTH_1(4,13));
			ADD_DEPTH_2(2,14)<=signed(ADD_DEPTH_1(3,14)) + signed(ADD_DEPTH_1(4,14));
			ADD_DEPTH_2(2,15)<=signed(ADD_DEPTH_1(3,15)) + signed(ADD_DEPTH_1(4,15));

			ADD_DEPTH_2(3,0)<=signed(ADD_DEPTH_1(5,0)) + signed(ADD_DEPTH_1(6,0));
			ADD_DEPTH_2(3,1)<=signed(ADD_DEPTH_1(5,1)) + signed(ADD_DEPTH_1(6,1));
			ADD_DEPTH_2(3,2)<=signed(ADD_DEPTH_1(5,2)) + signed(ADD_DEPTH_1(6,2));
			ADD_DEPTH_2(3,3)<=signed(ADD_DEPTH_1(5,3)) + signed(ADD_DEPTH_1(6,3));
			ADD_DEPTH_2(3,4)<=signed(ADD_DEPTH_1(5,4)) + signed(ADD_DEPTH_1(6,4));
			ADD_DEPTH_2(3,5)<=signed(ADD_DEPTH_1(5,5)) + signed(ADD_DEPTH_1(6,5));
			ADD_DEPTH_2(3,6)<=signed(ADD_DEPTH_1(5,6)) + signed(ADD_DEPTH_1(6,6));
			ADD_DEPTH_2(3,7)<=signed(ADD_DEPTH_1(5,7)) + signed(ADD_DEPTH_1(6,7));
			ADD_DEPTH_2(3,8)<=signed(ADD_DEPTH_1(5,8)) + signed(ADD_DEPTH_1(6,8));
			ADD_DEPTH_2(3,9)<=signed(ADD_DEPTH_1(5,9)) + signed(ADD_DEPTH_1(6,9));
			ADD_DEPTH_2(3,10)<=signed(ADD_DEPTH_1(5,10)) + signed(ADD_DEPTH_1(6,10));
			ADD_DEPTH_2(3,11)<=signed(ADD_DEPTH_1(5,11)) + signed(ADD_DEPTH_1(6,11));
			ADD_DEPTH_2(3,12)<=signed(ADD_DEPTH_1(5,12)) + signed(ADD_DEPTH_1(6,12));
			ADD_DEPTH_2(3,13)<=signed(ADD_DEPTH_1(5,13)) + signed(ADD_DEPTH_1(6,13));
			ADD_DEPTH_2(3,14)<=signed(ADD_DEPTH_1(5,14)) + signed(ADD_DEPTH_1(6,14));
			ADD_DEPTH_2(3,15)<=signed(ADD_DEPTH_1(5,15)) + signed(ADD_DEPTH_1(6,15));

			ADD_DEPTH_2(4,0)<=signed(ADD_DEPTH_1(7,0)) + signed(ADD_DEPTH_1(8,0));
			ADD_DEPTH_2(4,1)<=signed(ADD_DEPTH_1(7,1)) + signed(ADD_DEPTH_1(8,1));
			ADD_DEPTH_2(4,2)<=signed(ADD_DEPTH_1(7,2)) + signed(ADD_DEPTH_1(8,2));
			ADD_DEPTH_2(4,3)<=signed(ADD_DEPTH_1(7,3)) + signed(ADD_DEPTH_1(8,3));
			ADD_DEPTH_2(4,4)<=signed(ADD_DEPTH_1(7,4)) + signed(ADD_DEPTH_1(8,4));
			ADD_DEPTH_2(4,5)<=signed(ADD_DEPTH_1(7,5)) + signed(ADD_DEPTH_1(8,5));
			ADD_DEPTH_2(4,6)<=signed(ADD_DEPTH_1(7,6)) + signed(ADD_DEPTH_1(8,6));
			ADD_DEPTH_2(4,7)<=signed(ADD_DEPTH_1(7,7)) + signed(ADD_DEPTH_1(8,7));
			ADD_DEPTH_2(4,8)<=signed(ADD_DEPTH_1(7,8)) + signed(ADD_DEPTH_1(8,8));
			ADD_DEPTH_2(4,9)<=signed(ADD_DEPTH_1(7,9)) + signed(ADD_DEPTH_1(8,9));
			ADD_DEPTH_2(4,10)<=signed(ADD_DEPTH_1(7,10)) + signed(ADD_DEPTH_1(8,10));
			ADD_DEPTH_2(4,11)<=signed(ADD_DEPTH_1(7,11)) + signed(ADD_DEPTH_1(8,11));
			ADD_DEPTH_2(4,12)<=signed(ADD_DEPTH_1(7,12)) + signed(ADD_DEPTH_1(8,12));
			ADD_DEPTH_2(4,13)<=signed(ADD_DEPTH_1(7,13)) + signed(ADD_DEPTH_1(8,13));
			ADD_DEPTH_2(4,14)<=signed(ADD_DEPTH_1(7,14)) + signed(ADD_DEPTH_1(8,14));
			ADD_DEPTH_2(4,15)<=signed(ADD_DEPTH_1(7,15)) + signed(ADD_DEPTH_1(8,15));

			ADD_DEPTH_2(5,0)<=signed(ADD_DEPTH_1(9,0)) + signed(ADD_DEPTH_1(10,0));
			ADD_DEPTH_2(5,1)<=signed(ADD_DEPTH_1(9,1)) + signed(ADD_DEPTH_1(10,1));
			ADD_DEPTH_2(5,2)<=signed(ADD_DEPTH_1(9,2)) + signed(ADD_DEPTH_1(10,2));
			ADD_DEPTH_2(5,3)<=signed(ADD_DEPTH_1(9,3)) + signed(ADD_DEPTH_1(10,3));
			ADD_DEPTH_2(5,4)<=signed(ADD_DEPTH_1(9,4)) + signed(ADD_DEPTH_1(10,4));
			ADD_DEPTH_2(5,5)<=signed(ADD_DEPTH_1(9,5)) + signed(ADD_DEPTH_1(10,5));
			ADD_DEPTH_2(5,6)<=signed(ADD_DEPTH_1(9,6)) + signed(ADD_DEPTH_1(10,6));
			ADD_DEPTH_2(5,7)<=signed(ADD_DEPTH_1(9,7)) + signed(ADD_DEPTH_1(10,7));
			ADD_DEPTH_2(5,8)<=signed(ADD_DEPTH_1(9,8)) + signed(ADD_DEPTH_1(10,8));
			ADD_DEPTH_2(5,9)<=signed(ADD_DEPTH_1(9,9)) + signed(ADD_DEPTH_1(10,9));
			ADD_DEPTH_2(5,10)<=signed(ADD_DEPTH_1(9,10)) + signed(ADD_DEPTH_1(10,10));
			ADD_DEPTH_2(5,11)<=signed(ADD_DEPTH_1(9,11)) + signed(ADD_DEPTH_1(10,11));
			ADD_DEPTH_2(5,12)<=signed(ADD_DEPTH_1(9,12)) + signed(ADD_DEPTH_1(10,12));
			ADD_DEPTH_2(5,13)<=signed(ADD_DEPTH_1(9,13)) + signed(ADD_DEPTH_1(10,13));
			ADD_DEPTH_2(5,14)<=signed(ADD_DEPTH_1(9,14)) + signed(ADD_DEPTH_1(10,14));
			ADD_DEPTH_2(5,15)<=signed(ADD_DEPTH_1(9,15)) + signed(ADD_DEPTH_1(10,15));

			ADD_DEPTH_2(6,0)<=signed(ADD_DEPTH_1(11,0)) + signed(ADD_DEPTH_1(12,0));
			ADD_DEPTH_2(6,1)<=signed(ADD_DEPTH_1(11,1)) + signed(ADD_DEPTH_1(12,1));
			ADD_DEPTH_2(6,2)<=signed(ADD_DEPTH_1(11,2)) + signed(ADD_DEPTH_1(12,2));
			ADD_DEPTH_2(6,3)<=signed(ADD_DEPTH_1(11,3)) + signed(ADD_DEPTH_1(12,3));
			ADD_DEPTH_2(6,4)<=signed(ADD_DEPTH_1(11,4)) + signed(ADD_DEPTH_1(12,4));
			ADD_DEPTH_2(6,5)<=signed(ADD_DEPTH_1(11,5)) + signed(ADD_DEPTH_1(12,5));
			ADD_DEPTH_2(6,6)<=signed(ADD_DEPTH_1(11,6)) + signed(ADD_DEPTH_1(12,6));
			ADD_DEPTH_2(6,7)<=signed(ADD_DEPTH_1(11,7)) + signed(ADD_DEPTH_1(12,7));
			ADD_DEPTH_2(6,8)<=signed(ADD_DEPTH_1(11,8)) + signed(ADD_DEPTH_1(12,8));
			ADD_DEPTH_2(6,9)<=signed(ADD_DEPTH_1(11,9)) + signed(ADD_DEPTH_1(12,9));
			ADD_DEPTH_2(6,10)<=signed(ADD_DEPTH_1(11,10)) + signed(ADD_DEPTH_1(12,10));
			ADD_DEPTH_2(6,11)<=signed(ADD_DEPTH_1(11,11)) + signed(ADD_DEPTH_1(12,11));
			ADD_DEPTH_2(6,12)<=signed(ADD_DEPTH_1(11,12)) + signed(ADD_DEPTH_1(12,12));
			ADD_DEPTH_2(6,13)<=signed(ADD_DEPTH_1(11,13)) + signed(ADD_DEPTH_1(12,13));
			ADD_DEPTH_2(6,14)<=signed(ADD_DEPTH_1(11,14)) + signed(ADD_DEPTH_1(12,14));
			ADD_DEPTH_2(6,15)<=signed(ADD_DEPTH_1(11,15)) + signed(ADD_DEPTH_1(12,15));


				Enable_STAGE_3<= '1';
			end if; 
			------------------------------------STAGE-3--------------------------------------
		if Enable_STAGE_3 = '1' then

			ADD_DEPTH_3(0,0)<=signed(ADD_DEPTH_2(0,0));
			ADD_DEPTH_3(0,1)<=signed(ADD_DEPTH_2(0,1));
			ADD_DEPTH_3(0,2)<=signed(ADD_DEPTH_2(0,2));
			ADD_DEPTH_3(0,3)<=signed(ADD_DEPTH_2(0,3));
			ADD_DEPTH_3(0,4)<=signed(ADD_DEPTH_2(0,4));
			ADD_DEPTH_3(0,5)<=signed(ADD_DEPTH_2(0,5));
			ADD_DEPTH_3(0,6)<=signed(ADD_DEPTH_2(0,6));
			ADD_DEPTH_3(0,7)<=signed(ADD_DEPTH_2(0,7));
			ADD_DEPTH_3(0,8)<=signed(ADD_DEPTH_2(0,8));
			ADD_DEPTH_3(0,9)<=signed(ADD_DEPTH_2(0,9));
			ADD_DEPTH_3(0,10)<=signed(ADD_DEPTH_2(0,10));
			ADD_DEPTH_3(0,11)<=signed(ADD_DEPTH_2(0,11));
			ADD_DEPTH_3(0,12)<=signed(ADD_DEPTH_2(0,12));
			ADD_DEPTH_3(0,13)<=signed(ADD_DEPTH_2(0,13));
			ADD_DEPTH_3(0,14)<=signed(ADD_DEPTH_2(0,14));
			ADD_DEPTH_3(0,15)<=signed(ADD_DEPTH_2(0,15));

			ADD_DEPTH_3(1,0)<=signed(ADD_DEPTH_2(1,0)) + signed(ADD_DEPTH_2(2,0));
			ADD_DEPTH_3(1,1)<=signed(ADD_DEPTH_2(1,1)) + signed(ADD_DEPTH_2(2,1));
			ADD_DEPTH_3(1,2)<=signed(ADD_DEPTH_2(1,2)) + signed(ADD_DEPTH_2(2,2));
			ADD_DEPTH_3(1,3)<=signed(ADD_DEPTH_2(1,3)) + signed(ADD_DEPTH_2(2,3));
			ADD_DEPTH_3(1,4)<=signed(ADD_DEPTH_2(1,4)) + signed(ADD_DEPTH_2(2,4));
			ADD_DEPTH_3(1,5)<=signed(ADD_DEPTH_2(1,5)) + signed(ADD_DEPTH_2(2,5));
			ADD_DEPTH_3(1,6)<=signed(ADD_DEPTH_2(1,6)) + signed(ADD_DEPTH_2(2,6));
			ADD_DEPTH_3(1,7)<=signed(ADD_DEPTH_2(1,7)) + signed(ADD_DEPTH_2(2,7));
			ADD_DEPTH_3(1,8)<=signed(ADD_DEPTH_2(1,8)) + signed(ADD_DEPTH_2(2,8));
			ADD_DEPTH_3(1,9)<=signed(ADD_DEPTH_2(1,9)) + signed(ADD_DEPTH_2(2,9));
			ADD_DEPTH_3(1,10)<=signed(ADD_DEPTH_2(1,10)) + signed(ADD_DEPTH_2(2,10));
			ADD_DEPTH_3(1,11)<=signed(ADD_DEPTH_2(1,11)) + signed(ADD_DEPTH_2(2,11));
			ADD_DEPTH_3(1,12)<=signed(ADD_DEPTH_2(1,12)) + signed(ADD_DEPTH_2(2,12));
			ADD_DEPTH_3(1,13)<=signed(ADD_DEPTH_2(1,13)) + signed(ADD_DEPTH_2(2,13));
			ADD_DEPTH_3(1,14)<=signed(ADD_DEPTH_2(1,14)) + signed(ADD_DEPTH_2(2,14));
			ADD_DEPTH_3(1,15)<=signed(ADD_DEPTH_2(1,15)) + signed(ADD_DEPTH_2(2,15));

			ADD_DEPTH_3(2,0)<=signed(ADD_DEPTH_2(3,0)) + signed(ADD_DEPTH_2(4,0));
			ADD_DEPTH_3(2,1)<=signed(ADD_DEPTH_2(3,1)) + signed(ADD_DEPTH_2(4,1));
			ADD_DEPTH_3(2,2)<=signed(ADD_DEPTH_2(3,2)) + signed(ADD_DEPTH_2(4,2));
			ADD_DEPTH_3(2,3)<=signed(ADD_DEPTH_2(3,3)) + signed(ADD_DEPTH_2(4,3));
			ADD_DEPTH_3(2,4)<=signed(ADD_DEPTH_2(3,4)) + signed(ADD_DEPTH_2(4,4));
			ADD_DEPTH_3(2,5)<=signed(ADD_DEPTH_2(3,5)) + signed(ADD_DEPTH_2(4,5));
			ADD_DEPTH_3(2,6)<=signed(ADD_DEPTH_2(3,6)) + signed(ADD_DEPTH_2(4,6));
			ADD_DEPTH_3(2,7)<=signed(ADD_DEPTH_2(3,7)) + signed(ADD_DEPTH_2(4,7));
			ADD_DEPTH_3(2,8)<=signed(ADD_DEPTH_2(3,8)) + signed(ADD_DEPTH_2(4,8));
			ADD_DEPTH_3(2,9)<=signed(ADD_DEPTH_2(3,9)) + signed(ADD_DEPTH_2(4,9));
			ADD_DEPTH_3(2,10)<=signed(ADD_DEPTH_2(3,10)) + signed(ADD_DEPTH_2(4,10));
			ADD_DEPTH_3(2,11)<=signed(ADD_DEPTH_2(3,11)) + signed(ADD_DEPTH_2(4,11));
			ADD_DEPTH_3(2,12)<=signed(ADD_DEPTH_2(3,12)) + signed(ADD_DEPTH_2(4,12));
			ADD_DEPTH_3(2,13)<=signed(ADD_DEPTH_2(3,13)) + signed(ADD_DEPTH_2(4,13));
			ADD_DEPTH_3(2,14)<=signed(ADD_DEPTH_2(3,14)) + signed(ADD_DEPTH_2(4,14));
			ADD_DEPTH_3(2,15)<=signed(ADD_DEPTH_2(3,15)) + signed(ADD_DEPTH_2(4,15));

			ADD_DEPTH_3(3,0)<=signed(ADD_DEPTH_2(5,0)) + signed(ADD_DEPTH_2(6,0));
			ADD_DEPTH_3(3,1)<=signed(ADD_DEPTH_2(5,1)) + signed(ADD_DEPTH_2(6,1));
			ADD_DEPTH_3(3,2)<=signed(ADD_DEPTH_2(5,2)) + signed(ADD_DEPTH_2(6,2));
			ADD_DEPTH_3(3,3)<=signed(ADD_DEPTH_2(5,3)) + signed(ADD_DEPTH_2(6,3));
			ADD_DEPTH_3(3,4)<=signed(ADD_DEPTH_2(5,4)) + signed(ADD_DEPTH_2(6,4));
			ADD_DEPTH_3(3,5)<=signed(ADD_DEPTH_2(5,5)) + signed(ADD_DEPTH_2(6,5));
			ADD_DEPTH_3(3,6)<=signed(ADD_DEPTH_2(5,6)) + signed(ADD_DEPTH_2(6,6));
			ADD_DEPTH_3(3,7)<=signed(ADD_DEPTH_2(5,7)) + signed(ADD_DEPTH_2(6,7));
			ADD_DEPTH_3(3,8)<=signed(ADD_DEPTH_2(5,8)) + signed(ADD_DEPTH_2(6,8));
			ADD_DEPTH_3(3,9)<=signed(ADD_DEPTH_2(5,9)) + signed(ADD_DEPTH_2(6,9));
			ADD_DEPTH_3(3,10)<=signed(ADD_DEPTH_2(5,10)) + signed(ADD_DEPTH_2(6,10));
			ADD_DEPTH_3(3,11)<=signed(ADD_DEPTH_2(5,11)) + signed(ADD_DEPTH_2(6,11));
			ADD_DEPTH_3(3,12)<=signed(ADD_DEPTH_2(5,12)) + signed(ADD_DEPTH_2(6,12));
			ADD_DEPTH_3(3,13)<=signed(ADD_DEPTH_2(5,13)) + signed(ADD_DEPTH_2(6,13));
			ADD_DEPTH_3(3,14)<=signed(ADD_DEPTH_2(5,14)) + signed(ADD_DEPTH_2(6,14));
			ADD_DEPTH_3(3,15)<=signed(ADD_DEPTH_2(5,15)) + signed(ADD_DEPTH_2(6,15));


				Enable_STAGE_4<= '1';
			end if; 
			------------------------------------STAGE-4--------------------------------------
		if Enable_STAGE_4 = '1' then


			ADD_DEPTH_4(0,0)<=signed(ADD_DEPTH_3(0,0)) + signed(ADD_DEPTH_3(1,0));
			ADD_DEPTH_4(0,1)<=signed(ADD_DEPTH_3(0,1)) + signed(ADD_DEPTH_3(1,1));
			ADD_DEPTH_4(0,2)<=signed(ADD_DEPTH_3(0,2)) + signed(ADD_DEPTH_3(1,2));
			ADD_DEPTH_4(0,3)<=signed(ADD_DEPTH_3(0,3)) + signed(ADD_DEPTH_3(1,3));
			ADD_DEPTH_4(0,4)<=signed(ADD_DEPTH_3(0,4)) + signed(ADD_DEPTH_3(1,4));
			ADD_DEPTH_4(0,5)<=signed(ADD_DEPTH_3(0,5)) + signed(ADD_DEPTH_3(1,5));
			ADD_DEPTH_4(0,6)<=signed(ADD_DEPTH_3(0,6)) + signed(ADD_DEPTH_3(1,6));
			ADD_DEPTH_4(0,7)<=signed(ADD_DEPTH_3(0,7)) + signed(ADD_DEPTH_3(1,7));
			ADD_DEPTH_4(0,8)<=signed(ADD_DEPTH_3(0,8)) + signed(ADD_DEPTH_3(1,8));
			ADD_DEPTH_4(0,9)<=signed(ADD_DEPTH_3(0,9)) + signed(ADD_DEPTH_3(1,9));
			ADD_DEPTH_4(0,10)<=signed(ADD_DEPTH_3(0,10)) + signed(ADD_DEPTH_3(1,10));
			ADD_DEPTH_4(0,11)<=signed(ADD_DEPTH_3(0,11)) + signed(ADD_DEPTH_3(1,11));
			ADD_DEPTH_4(0,12)<=signed(ADD_DEPTH_3(0,12)) + signed(ADD_DEPTH_3(1,12));
			ADD_DEPTH_4(0,13)<=signed(ADD_DEPTH_3(0,13)) + signed(ADD_DEPTH_3(1,13));
			ADD_DEPTH_4(0,14)<=signed(ADD_DEPTH_3(0,14)) + signed(ADD_DEPTH_3(1,14));
			ADD_DEPTH_4(0,15)<=signed(ADD_DEPTH_3(0,15)) + signed(ADD_DEPTH_3(1,15));

			ADD_DEPTH_4(1,0)<=signed(ADD_DEPTH_3(2,0)) + signed(ADD_DEPTH_3(3,0));
			ADD_DEPTH_4(1,1)<=signed(ADD_DEPTH_3(2,1)) + signed(ADD_DEPTH_3(3,1));
			ADD_DEPTH_4(1,2)<=signed(ADD_DEPTH_3(2,2)) + signed(ADD_DEPTH_3(3,2));
			ADD_DEPTH_4(1,3)<=signed(ADD_DEPTH_3(2,3)) + signed(ADD_DEPTH_3(3,3));
			ADD_DEPTH_4(1,4)<=signed(ADD_DEPTH_3(2,4)) + signed(ADD_DEPTH_3(3,4));
			ADD_DEPTH_4(1,5)<=signed(ADD_DEPTH_3(2,5)) + signed(ADD_DEPTH_3(3,5));
			ADD_DEPTH_4(1,6)<=signed(ADD_DEPTH_3(2,6)) + signed(ADD_DEPTH_3(3,6));
			ADD_DEPTH_4(1,7)<=signed(ADD_DEPTH_3(2,7)) + signed(ADD_DEPTH_3(3,7));
			ADD_DEPTH_4(1,8)<=signed(ADD_DEPTH_3(2,8)) + signed(ADD_DEPTH_3(3,8));
			ADD_DEPTH_4(1,9)<=signed(ADD_DEPTH_3(2,9)) + signed(ADD_DEPTH_3(3,9));
			ADD_DEPTH_4(1,10)<=signed(ADD_DEPTH_3(2,10)) + signed(ADD_DEPTH_3(3,10));
			ADD_DEPTH_4(1,11)<=signed(ADD_DEPTH_3(2,11)) + signed(ADD_DEPTH_3(3,11));
			ADD_DEPTH_4(1,12)<=signed(ADD_DEPTH_3(2,12)) + signed(ADD_DEPTH_3(3,12));
			ADD_DEPTH_4(1,13)<=signed(ADD_DEPTH_3(2,13)) + signed(ADD_DEPTH_3(3,13));
			ADD_DEPTH_4(1,14)<=signed(ADD_DEPTH_3(2,14)) + signed(ADD_DEPTH_3(3,14));
			ADD_DEPTH_4(1,15)<=signed(ADD_DEPTH_3(2,15)) + signed(ADD_DEPTH_3(3,15));


				Enable_STAGE_5<= '1';
			end if; 
			------------------------------------STAGE-5--------------------------------------
		if Enable_STAGE_5 = '1' then


			ADD_DEPTH_5(0,0)<=signed(ADD_DEPTH_4(0,0)) + signed(ADD_DEPTH_4(1,0));
			ADD_DEPTH_5(0,1)<=signed(ADD_DEPTH_4(0,1)) + signed(ADD_DEPTH_4(1,1));
			ADD_DEPTH_5(0,2)<=signed(ADD_DEPTH_4(0,2)) + signed(ADD_DEPTH_4(1,2));
			ADD_DEPTH_5(0,3)<=signed(ADD_DEPTH_4(0,3)) + signed(ADD_DEPTH_4(1,3));
			ADD_DEPTH_5(0,4)<=signed(ADD_DEPTH_4(0,4)) + signed(ADD_DEPTH_4(1,4));
			ADD_DEPTH_5(0,5)<=signed(ADD_DEPTH_4(0,5)) + signed(ADD_DEPTH_4(1,5));
			ADD_DEPTH_5(0,6)<=signed(ADD_DEPTH_4(0,6)) + signed(ADD_DEPTH_4(1,6));
			ADD_DEPTH_5(0,7)<=signed(ADD_DEPTH_4(0,7)) + signed(ADD_DEPTH_4(1,7));
			ADD_DEPTH_5(0,8)<=signed(ADD_DEPTH_4(0,8)) + signed(ADD_DEPTH_4(1,8));
			ADD_DEPTH_5(0,9)<=signed(ADD_DEPTH_4(0,9)) + signed(ADD_DEPTH_4(1,9));
			ADD_DEPTH_5(0,10)<=signed(ADD_DEPTH_4(0,10)) + signed(ADD_DEPTH_4(1,10));
			ADD_DEPTH_5(0,11)<=signed(ADD_DEPTH_4(0,11)) + signed(ADD_DEPTH_4(1,11));
			ADD_DEPTH_5(0,12)<=signed(ADD_DEPTH_4(0,12)) + signed(ADD_DEPTH_4(1,12));
			ADD_DEPTH_5(0,13)<=signed(ADD_DEPTH_4(0,13)) + signed(ADD_DEPTH_4(1,13));
			ADD_DEPTH_5(0,14)<=signed(ADD_DEPTH_4(0,14)) + signed(ADD_DEPTH_4(1,14));
			ADD_DEPTH_5(0,15)<=signed(ADD_DEPTH_4(0,15)) + signed(ADD_DEPTH_4(1,15));


			Enable_BIAS<='1'; 
		end if;
		------------------------------------STAGE-BIAS--------------------------------------
		
		if Enable_BIAS = '1' then

			BIAS_1<=(signed(BIAS_VAL_1)+signed(ADD_DEPTH_5(0,0)(PERCISION downto 1)));
			BIAS_2<=(signed(BIAS_VAL_2)+signed(ADD_DEPTH_5(0,1)(PERCISION downto 1)));
			BIAS_3<=(signed(BIAS_VAL_3)+signed(ADD_DEPTH_5(0,2)(PERCISION downto 1)));
			BIAS_4<=(signed(BIAS_VAL_4)+signed(ADD_DEPTH_5(0,3)(PERCISION downto 1)));
			BIAS_5<=(signed(BIAS_VAL_5)+signed(ADD_DEPTH_5(0,4)(PERCISION downto 1)));
			BIAS_6<=(signed(BIAS_VAL_6)+signed(ADD_DEPTH_5(0,5)(PERCISION downto 1)));
			BIAS_7<=(signed(BIAS_VAL_7)+signed(ADD_DEPTH_5(0,6)(PERCISION downto 1)));
			BIAS_8<=(signed(BIAS_VAL_8)+signed(ADD_DEPTH_5(0,7)(PERCISION downto 1)));
			BIAS_9<=(signed(BIAS_VAL_9)+signed(ADD_DEPTH_5(0,8)(PERCISION downto 1)));
			BIAS_10<=(signed(BIAS_VAL_10)+signed(ADD_DEPTH_5(0,9)(PERCISION downto 1)));
			BIAS_11<=(signed(BIAS_VAL_11)+signed(ADD_DEPTH_5(0,10)(PERCISION downto 1)));
			BIAS_12<=(signed(BIAS_VAL_12)+signed(ADD_DEPTH_5(0,11)(PERCISION downto 1)));
			BIAS_13<=(signed(BIAS_VAL_13)+signed(ADD_DEPTH_5(0,12)(PERCISION downto 1)));
			BIAS_14<=(signed(BIAS_VAL_14)+signed(ADD_DEPTH_5(0,13)(PERCISION downto 1)));
			BIAS_15<=(signed(BIAS_VAL_15)+signed(ADD_DEPTH_5(0,14)(PERCISION downto 1)));
			BIAS_16<=(signed(BIAS_VAL_16)+signed(ADD_DEPTH_5(0,15)(PERCISION downto 1)));

			Enable_ReLU<='1';
			
		end if;

		if SIG_STRIDE>1 and Enable_ReLU='1' then
                 SIG_STRIDE<=SIG_STRIDE-1;
               elsif VALID_NXTLYR_PIX<(IMAGE_WIDTH-F_SIZE) then
		 SIG_STRIDE<=STRIDE; end if;

	if  Enable_ReLU='1' then
		if SIG_STRIDE>(STRIDE-1) and VALID_NXTLYR_PIX<=(IMAGE_WIDTH-F_SIZE) then          --VALID_NXTLYR_PIX<IMAGE_WIDTH and  VALID_LOCAL_PIX

			if BIAS_1>0 then
			ReLU_1<=BIAS_1;
			DOUT_BUF_1_3<=std_logic_vector(BIAS_1);
			else
			ReLU_1<= (others => '0');
			DOUT_BUF_1_3<=(others => '0');
			end if;
			if BIAS_2>0 then
			ReLU_2<=BIAS_2;
			DOUT_BUF_2_3<=std_logic_vector(BIAS_2);
			else
			ReLU_2<= (others => '0');
			DOUT_BUF_2_3<=(others => '0');
			end if;
			if BIAS_3>0 then
			ReLU_3<=BIAS_3;
			DOUT_BUF_3_3<=std_logic_vector(BIAS_3);
			else
			ReLU_3<= (others => '0');
			DOUT_BUF_3_3<=(others => '0');
			end if;
			if BIAS_4>0 then
			ReLU_4<=BIAS_4;
			DOUT_BUF_4_3<=std_logic_vector(BIAS_4);
			else
			ReLU_4<= (others => '0');
			DOUT_BUF_4_3<=(others => '0');
			end if;
			if BIAS_5>0 then
			ReLU_5<=BIAS_5;
			DOUT_BUF_5_3<=std_logic_vector(BIAS_5);
			else
			ReLU_5<= (others => '0');
			DOUT_BUF_5_3<=(others => '0');
			end if;
			if BIAS_6>0 then
			ReLU_6<=BIAS_6;
			DOUT_BUF_6_3<=std_logic_vector(BIAS_6);
			else
			ReLU_6<= (others => '0');
			DOUT_BUF_6_3<=(others => '0');
			end if;
			if BIAS_7>0 then
			ReLU_7<=BIAS_7;
			DOUT_BUF_7_3<=std_logic_vector(BIAS_7);
			else
			ReLU_7<= (others => '0');
			DOUT_BUF_7_3<=(others => '0');
			end if;
			if BIAS_8>0 then
			ReLU_8<=BIAS_8;
			DOUT_BUF_8_3<=std_logic_vector(BIAS_8);
			else
			ReLU_8<= (others => '0');
			DOUT_BUF_8_3<=(others => '0');
			end if;
			if BIAS_9>0 then
			ReLU_9<=BIAS_9;
			DOUT_BUF_9_3<=std_logic_vector(BIAS_9);
			else
			ReLU_9<= (others => '0');
			DOUT_BUF_9_3<=(others => '0');
			end if;
			if BIAS_10>0 then
			ReLU_10<=BIAS_10;
			DOUT_BUF_10_3<=std_logic_vector(BIAS_10);
			else
			ReLU_10<= (others => '0');
			DOUT_BUF_10_3<=(others => '0');
			end if;
			if BIAS_11>0 then
			ReLU_11<=BIAS_11;
			DOUT_BUF_11_3<=std_logic_vector(BIAS_11);
			else
			ReLU_11<= (others => '0');
			DOUT_BUF_11_3<=(others => '0');
			end if;
			if BIAS_12>0 then
			ReLU_12<=BIAS_12;
			DOUT_BUF_12_3<=std_logic_vector(BIAS_12);
			else
			ReLU_12<= (others => '0');
			DOUT_BUF_12_3<=(others => '0');
			end if;
			if BIAS_13>0 then
			ReLU_13<=BIAS_13;
			DOUT_BUF_13_3<=std_logic_vector(BIAS_13);
			else
			ReLU_13<= (others => '0');
			DOUT_BUF_13_3<=(others => '0');
			end if;
			if BIAS_14>0 then
			ReLU_14<=BIAS_14;
			DOUT_BUF_14_3<=std_logic_vector(BIAS_14);
			else
			ReLU_14<= (others => '0');
			DOUT_BUF_14_3<=(others => '0');
			end if;
			if BIAS_15>0 then
			ReLU_15<=BIAS_15;
			DOUT_BUF_15_3<=std_logic_vector(BIAS_15);
			else
			ReLU_15<= (others => '0');
			DOUT_BUF_15_3<=(others => '0');
			end if;
			if BIAS_16>0 then
			ReLU_16<=BIAS_16;
			DOUT_BUF_16_3<=std_logic_vector(BIAS_16);
			else
			ReLU_16<= (others => '0');
			DOUT_BUF_16_3<=(others => '0');
			end if;

			EN_NXT_LYR_3<='1';FRST_TIM_EN_3<='1';
			OUT_PIXEL_COUNT<=OUT_PIXEL_COUNT+1;
		else
               EN_NXT_LYR_3<='0';
               DOUT_BUF_1_3<=(others => '0');
               DOUT_BUF_2_3<=(others => '0');
               DOUT_BUF_3_3<=(others => '0');
               DOUT_BUF_4_3<=(others => '0');
               DOUT_BUF_5_3<=(others => '0');
               DOUT_BUF_6_3<=(others => '0');
               DOUT_BUF_7_3<=(others => '0');
               DOUT_BUF_8_3<=(others => '0');
               DOUT_BUF_9_3<=(others => '0');
               DOUT_BUF_10_3<=(others => '0');
               DOUT_BUF_11_3<=(others => '0');
               DOUT_BUF_12_3<=(others => '0');
               DOUT_BUF_13_3<=(others => '0');
               DOUT_BUF_14_3<=(others => '0');
               DOUT_BUF_15_3<=(others => '0');
               DOUT_BUF_16_3<=(others => '0');

		end if; -- VALIDPIXELS

		if VALID_NXTLYR_PIX=((IMAGE_WIDTH*STRIDE)-1) then VALID_NXTLYR_PIX<=0;SIG_STRIDE<=STRIDE;   -- reset sride and valid pixels
		else VALID_NXTLYR_PIX<=VALID_NXTLYR_PIX+1;end if; 

	end if;  --ReLU

	--end if;  --enable window              canceled 

 elsif OUT_PIXEL_COUNT>=VALID_CYCLES  then INTERNAL_RST<='1';SIG_STRIDE<=STRIDE;EN_NXT_LYR_3<='1';  -- order is very important
else  EN_NXT_LYR_3<='0';-- In case stream stopped

end if; -- end enable 
end if; -- for RST	
end if; -- rising edge
end process LAYER_3;

EN_STREAM_OUT_3<= EN_STREAM_OUT_4;
VALID_OUT_3<= VALID_OUT_4;
DOUT_1_3<=DOUT_1_4;
DOUT_2_3<=DOUT_2_4;
DOUT_3_3<=DOUT_3_4;
DOUT_4_3<=DOUT_4_4;
DOUT_5_3<=DOUT_5_4;
DOUT_6_3<=DOUT_6_4;
DOUT_7_3<=DOUT_7_4;
DOUT_8_3<=DOUT_8_4;
DOUT_9_3<=DOUT_9_4;
DOUT_10_3<=DOUT_10_4;

end Behavioral;
------------------------------ ARCHITECTURE DECLARATION - END---------------------------------------------

